module GunzipBitSkipper( // @[:@3.2]
  input   clock, // @[:@4.4]
  input   reset, // @[:@5.4]
  input   io_data_in_valid, // @[:@6.4]
  output  io_data_in_ready, // @[:@6.4]
  output  io_done // @[:@6.4]
);
  reg [8:0] bit_cntr; // @[GunzipBitSkipper.scala 43:25:@8.4]
  reg [31:0] _RAND_0;
  wire  _T_13; // @[GunzipBitSkipper.scala 45:26:@9.4]
  wire  _T_15; // @[GunzipBitSkipper.scala 45:58:@10.4]
  wire  _T_16; // @[GunzipBitSkipper.scala 45:46:@11.4]
  wire [9:0] _T_18; // @[GunzipBitSkipper.scala 46:26:@13.6]
  wire [8:0] _T_19; // @[GunzipBitSkipper.scala 46:26:@14.6]
  wire [8:0] _GEN_0; // @[GunzipBitSkipper.scala 45:80:@12.4]
  assign _T_13 = io_data_in_ready & io_data_in_valid; // @[GunzipBitSkipper.scala 45:26:@9.4]
  assign _T_15 = bit_cntr < 9'h1a7; // @[GunzipBitSkipper.scala 45:58:@10.4]
  assign _T_16 = _T_13 & _T_15; // @[GunzipBitSkipper.scala 45:46:@11.4]
  assign _T_18 = bit_cntr + 9'h1; // @[GunzipBitSkipper.scala 46:26:@13.6]
  assign _T_19 = bit_cntr + 9'h1; // @[GunzipBitSkipper.scala 46:26:@14.6]
  assign _GEN_0 = _T_16 ? _T_19 : bit_cntr; // @[GunzipBitSkipper.scala 45:80:@12.4]
  assign io_data_in_ready = bit_cntr != 9'h1a7; // @[GunzipBitSkipper.scala 50:20:@20.4]
  assign io_done = bit_cntr == 9'h1a7; // @[GunzipBitSkipper.scala 49:11:@18.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bit_cntr = _RAND_0[8:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      bit_cntr <= 9'h0;
    end else begin
      if (_T_16) begin
        bit_cntr <= _T_19;
      end
    end
  end
endmodule
module GunzipHuffDecoder( // @[:@22.2]
  input        clock, // @[:@23.4]
  input        reset, // @[:@24.4]
  input        io_data_in_valid, // @[:@25.4]
  output       io_data_in_ready, // @[:@25.4]
  input        io_data_in_bits, // @[:@25.4]
  input        io_enable, // @[:@25.4]
  output [8:0] io_data, // @[:@25.4]
  output       io_valid // @[:@25.4]
);
  reg [8:0] lit_idx; // @[GunzipHuffDecoder.scala 41:24:@27.4]
  reg [31:0] _RAND_0;
  reg [8:0] data_reg; // @[GunzipHuffDecoder.scala 43:21:@539.4]
  reg [31:0] _RAND_1;
  wire  _T_794; // @[GunzipHuffDecoder.scala 52:19:@546.6]
  wire  _T_797; // @[GunzipHuffDecoder.scala 54:13:@549.8]
  wire [10:0] _T_800; // @[GunzipHuffDecoder.scala 58:25:@557.10]
  wire [11:0] _T_802; // @[GunzipHuffDecoder.scala 58:30:@558.10]
  wire [10:0] _T_803; // @[GunzipHuffDecoder.scala 58:30:@559.10]
  wire [10:0] _GEN_1550; // @[GunzipHuffDecoder.scala 58:36:@560.10]
  wire [11:0] _T_804; // @[GunzipHuffDecoder.scala 58:36:@560.10]
  wire [10:0] _T_805; // @[GunzipHuffDecoder.scala 58:36:@561.10]
  wire [7:0] _T_807; // @[:@563.10]
  wire  _GEN_6; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_7; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_8; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_9; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_10; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_11; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_12; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_13; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_14; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_15; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_16; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_17; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_18; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_19; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_20; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_21; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_22; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_23; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_24; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_25; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_26; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_27; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_28; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_29; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_30; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_31; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_32; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_33; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_34; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_35; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_36; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_37; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_38; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_39; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_40; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_41; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_42; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_43; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_44; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_45; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_46; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_47; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_48; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_49; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_50; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_51; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_52; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_53; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_54; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_55; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_56; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_57; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_58; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_59; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_60; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_61; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_62; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_63; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_64; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_65; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_66; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_67; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_68; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_69; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_70; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_71; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_72; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_73; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_74; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_75; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_76; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_77; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_78; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_79; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_80; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_81; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_82; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_83; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_84; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_85; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_86; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_87; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_88; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_89; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_90; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_91; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_92; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_93; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_94; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_95; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_96; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_97; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_98; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_99; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_100; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_101; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_102; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_103; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_104; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_105; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_106; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_107; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_108; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_109; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_110; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_111; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_112; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_113; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_114; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_115; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_116; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_117; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_118; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_119; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_120; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_121; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_122; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_123; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_124; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_125; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_126; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_127; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_128; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_129; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_130; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_131; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_132; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_133; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_134; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_135; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_136; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_137; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_138; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_139; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_140; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_141; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_142; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_143; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_144; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_145; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_146; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_147; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_148; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_149; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_150; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_151; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_152; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_153; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_154; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_155; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_156; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_157; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_158; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_159; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_160; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_161; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_162; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_163; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_164; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_165; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_166; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_167; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_168; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_169; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_170; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_171; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_172; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_173; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_174; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_175; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_176; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_177; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_178; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_179; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_180; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_181; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_182; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_183; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_184; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_185; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_186; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_187; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_188; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_189; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_190; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_191; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_192; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_193; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_194; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_195; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_196; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_197; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_198; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_199; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_200; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_201; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_202; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_203; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_204; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_205; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_206; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_207; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_208; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_209; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_210; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_211; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_212; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_213; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_214; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_215; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_216; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_217; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_218; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_219; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_220; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_221; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_222; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_223; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_224; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_225; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_226; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_227; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_228; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_229; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_230; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_231; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_232; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_233; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_234; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_235; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_236; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_237; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_238; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_239; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_240; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_241; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_242; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_243; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_244; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_245; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_246; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_247; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_248; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_249; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_250; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_251; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_252; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_253; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_254; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_255; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_256; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_257; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_258; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_259; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_260; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_261; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_262; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_263; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_264; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_265; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_266; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_267; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_268; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_269; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_270; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_271; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_272; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_273; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_274; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_275; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_276; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_277; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_278; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_279; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_280; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_281; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_282; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_283; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_284; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_285; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_286; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_287; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_288; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_289; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_290; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_291; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_292; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_293; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_294; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_295; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_296; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_297; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_298; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_299; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_300; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_301; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_302; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_303; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_304; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_305; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_306; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_307; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_308; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_309; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_310; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_311; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_312; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_313; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_314; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_315; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_316; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_317; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_318; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_319; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_320; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_321; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_322; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_323; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_324; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_325; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_326; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_327; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_328; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_329; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_330; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_331; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_332; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_333; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_334; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_335; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_336; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_337; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_338; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_339; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_340; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_341; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_342; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_343; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_344; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_345; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_346; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_347; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_348; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_349; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_350; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_351; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_352; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_353; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_354; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_355; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_356; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_357; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_358; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_359; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_360; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_361; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_362; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_363; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_364; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_365; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_366; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_367; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_368; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_369; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_370; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_371; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_372; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_373; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_374; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_375; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_376; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_377; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_378; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_379; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_380; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_381; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_382; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_383; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_384; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_385; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_386; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_387; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_388; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_389; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_390; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_391; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_392; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_393; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_394; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_395; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_396; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_397; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_398; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_399; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_400; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_401; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_402; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_403; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_404; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_405; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_406; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_407; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_408; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_409; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_410; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_411; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_412; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_413; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_414; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_415; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_416; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_417; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_418; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_419; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_420; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_421; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_422; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_423; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_424; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_425; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_426; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_427; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_428; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_429; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_430; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_431; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_432; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_433; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_434; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_435; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_436; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_437; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_438; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_439; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_440; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_441; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_442; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_443; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_444; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_445; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_446; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_447; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_448; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_449; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_450; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_451; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_452; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_453; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_454; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_455; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_456; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_457; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_458; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_459; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_460; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_461; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_462; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_463; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_464; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_465; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_466; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_467; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_468; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_469; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_470; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_471; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_472; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_473; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_474; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_475; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_476; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_477; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_478; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_479; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_480; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_481; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_482; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_483; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_484; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_485; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_486; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_487; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_488; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_489; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_490; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_491; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_492; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_493; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_494; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_495; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_496; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_497; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_498; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_499; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_500; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_501; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_502; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_503; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_504; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_505; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_506; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_507; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_508; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_509; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [10:0] _GEN_1530; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_1531; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire [8:0] _GEN_1532; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  wire  _GEN_1535; // @[GunzipHuffDecoder.scala 55:29:@555.8]
  wire [10:0] _GEN_1536; // @[GunzipHuffDecoder.scala 55:29:@555.8]
  wire [8:0] _GEN_1537; // @[GunzipHuffDecoder.scala 55:29:@555.8]
  wire  _GEN_1539; // @[GunzipHuffDecoder.scala 55:29:@555.8]
  wire  _GEN_1540; // @[GunzipHuffDecoder.scala 52:46:@547.6]
  wire [10:0] _GEN_1541; // @[GunzipHuffDecoder.scala 52:46:@547.6]
  wire [8:0] _GEN_1542; // @[GunzipHuffDecoder.scala 52:46:@547.6]
  wire  _GEN_1544; // @[GunzipHuffDecoder.scala 52:46:@547.6]
  wire [10:0] _GEN_1546; // @[GunzipHuffDecoder.scala 51:27:@545.4]
  wire  _GEN_1551; // @[GunzipHuffDecoder.scala 54:13:@551.10]
  assign _T_794 = lit_idx >= 9'hff; // @[GunzipHuffDecoder.scala 52:19:@546.6]
  assign _T_797 = reset == 1'h0; // @[GunzipHuffDecoder.scala 54:13:@549.8]
  assign _T_800 = lit_idx * 9'h2; // @[GunzipHuffDecoder.scala 58:25:@557.10]
  assign _T_802 = _T_800 + 11'h1; // @[GunzipHuffDecoder.scala 58:30:@558.10]
  assign _T_803 = _T_800 + 11'h1; // @[GunzipHuffDecoder.scala 58:30:@559.10]
  assign _GEN_1550 = {{10'd0}, io_data_in_bits}; // @[GunzipHuffDecoder.scala 58:36:@560.10]
  assign _T_804 = _T_803 + _GEN_1550; // @[GunzipHuffDecoder.scala 58:36:@560.10]
  assign _T_805 = _T_803 + _GEN_1550; // @[GunzipHuffDecoder.scala 58:36:@561.10]
  assign _T_807 = lit_idx[7:0]; // @[:@563.10]
  assign _GEN_6 = 8'h3 == _T_807; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_7 = 8'h3 == _T_807 ? 9'h11d : 9'h0; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_8 = 8'h4 == _T_807 ? 1'h0 : _GEN_6; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_9 = 8'h4 == _T_807 ? 9'h0 : _GEN_7; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_10 = 8'h5 == _T_807 ? 1'h0 : _GEN_8; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_11 = 8'h5 == _T_807 ? 9'h0 : _GEN_9; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_12 = 8'h6 == _T_807 ? 1'h0 : _GEN_10; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_13 = 8'h6 == _T_807 ? 9'h0 : _GEN_11; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_14 = 8'h7 == _T_807 ? 1'h0 : _GEN_12; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_15 = 8'h7 == _T_807 ? 9'h0 : _GEN_13; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_16 = 8'h8 == _T_807 ? 1'h0 : _GEN_14; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_17 = 8'h8 == _T_807 ? 9'h0 : _GEN_15; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_18 = 8'h9 == _T_807 ? 1'h0 : _GEN_16; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_19 = 8'h9 == _T_807 ? 9'h0 : _GEN_17; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_20 = 8'ha == _T_807 ? 1'h0 : _GEN_18; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_21 = 8'ha == _T_807 ? 9'h0 : _GEN_19; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_22 = 8'hb == _T_807 ? 1'h0 : _GEN_20; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_23 = 8'hb == _T_807 ? 9'h0 : _GEN_21; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_24 = 8'hc == _T_807 ? 1'h0 : _GEN_22; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_25 = 8'hc == _T_807 ? 9'h0 : _GEN_23; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_26 = 8'hd == _T_807 ? 1'h0 : _GEN_24; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_27 = 8'hd == _T_807 ? 9'h0 : _GEN_25; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_28 = 8'he == _T_807 ? 1'h0 : _GEN_26; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_29 = 8'he == _T_807 ? 9'h0 : _GEN_27; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_30 = 8'hf == _T_807 ? 1'h0 : _GEN_28; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_31 = 8'hf == _T_807 ? 9'h0 : _GEN_29; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_32 = 8'h10 == _T_807 ? 1'h0 : _GEN_30; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_33 = 8'h10 == _T_807 ? 9'h0 : _GEN_31; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_34 = 8'h11 == _T_807 ? 1'h0 : _GEN_32; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_35 = 8'h11 == _T_807 ? 9'h0 : _GEN_33; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_36 = 8'h12 == _T_807 ? 1'h0 : _GEN_34; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_37 = 8'h12 == _T_807 ? 9'h0 : _GEN_35; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_38 = 8'h13 == _T_807 ? 1'h1 : _GEN_36; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_39 = 8'h13 == _T_807 ? 9'h20 : _GEN_37; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_40 = 8'h14 == _T_807 ? 1'h1 : _GEN_38; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_41 = 8'h14 == _T_807 ? 9'h74 : _GEN_39; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_42 = 8'h15 == _T_807 ? 1'h0 : _GEN_40; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_43 = 8'h15 == _T_807 ? 9'h0 : _GEN_41; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_44 = 8'h16 == _T_807 ? 1'h0 : _GEN_42; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_45 = 8'h16 == _T_807 ? 9'h0 : _GEN_43; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_46 = 8'h17 == _T_807 ? 1'h0 : _GEN_44; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_47 = 8'h17 == _T_807 ? 9'h0 : _GEN_45; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_48 = 8'h18 == _T_807 ? 1'h0 : _GEN_46; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_49 = 8'h18 == _T_807 ? 9'h0 : _GEN_47; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_50 = 8'h19 == _T_807 ? 1'h0 : _GEN_48; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_51 = 8'h19 == _T_807 ? 9'h0 : _GEN_49; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_52 = 8'h1a == _T_807 ? 1'h0 : _GEN_50; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_53 = 8'h1a == _T_807 ? 9'h0 : _GEN_51; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_54 = 8'h1b == _T_807 ? 1'h0 : _GEN_52; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_55 = 8'h1b == _T_807 ? 9'h0 : _GEN_53; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_56 = 8'h1c == _T_807 ? 1'h0 : _GEN_54; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_57 = 8'h1c == _T_807 ? 9'h0 : _GEN_55; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_58 = 8'h1d == _T_807 ? 1'h0 : _GEN_56; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_59 = 8'h1d == _T_807 ? 9'h0 : _GEN_57; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_60 = 8'h1e == _T_807 ? 1'h0 : _GEN_58; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_61 = 8'h1e == _T_807 ? 9'h0 : _GEN_59; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_62 = 8'h1f == _T_807 ? 1'h0 : _GEN_60; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_63 = 8'h1f == _T_807 ? 9'h0 : _GEN_61; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_64 = 8'h20 == _T_807 ? 1'h0 : _GEN_62; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_65 = 8'h20 == _T_807 ? 9'h0 : _GEN_63; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_66 = 8'h21 == _T_807 ? 1'h0 : _GEN_64; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_67 = 8'h21 == _T_807 ? 9'h0 : _GEN_65; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_68 = 8'h22 == _T_807 ? 1'h0 : _GEN_66; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_69 = 8'h22 == _T_807 ? 9'h0 : _GEN_67; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_70 = 8'h23 == _T_807 ? 1'h0 : _GEN_68; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_71 = 8'h23 == _T_807 ? 9'h0 : _GEN_69; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_72 = 8'h24 == _T_807 ? 1'h0 : _GEN_70; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_73 = 8'h24 == _T_807 ? 9'h0 : _GEN_71; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_74 = 8'h25 == _T_807 ? 1'h0 : _GEN_72; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_75 = 8'h25 == _T_807 ? 9'h0 : _GEN_73; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_76 = 8'h26 == _T_807 ? 1'h0 : _GEN_74; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_77 = 8'h26 == _T_807 ? 9'h0 : _GEN_75; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_78 = 8'h27 == _T_807 ? 1'h0 : _GEN_76; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_79 = 8'h27 == _T_807 ? 9'h0 : _GEN_77; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_80 = 8'h28 == _T_807 ? 1'h0 : _GEN_78; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_81 = 8'h28 == _T_807 ? 9'h0 : _GEN_79; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_82 = 8'h29 == _T_807 ? 1'h0 : _GEN_80; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_83 = 8'h29 == _T_807 ? 9'h0 : _GEN_81; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_84 = 8'h2a == _T_807 ? 1'h0 : _GEN_82; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_85 = 8'h2a == _T_807 ? 9'h0 : _GEN_83; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_86 = 8'h2b == _T_807 ? 1'h1 : _GEN_84; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_87 = 8'h2b == _T_807 ? 9'h0 : _GEN_85; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_88 = 8'h2c == _T_807 ? 1'h1 : _GEN_86; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_89 = 8'h2c == _T_807 ? 9'ha : _GEN_87; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_90 = 8'h2d == _T_807 ? 1'h1 : _GEN_88; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_91 = 8'h2d == _T_807 ? 9'h31 : _GEN_89; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_92 = 8'h2e == _T_807 ? 1'h1 : _GEN_90; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_93 = 8'h2e == _T_807 ? 9'h33 : _GEN_91; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_94 = 8'h2f == _T_807 ? 1'h1 : _GEN_92; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_95 = 8'h2f == _T_807 ? 9'h34 : _GEN_93; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_96 = 8'h30 == _T_807 ? 1'h1 : _GEN_94; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_97 = 8'h30 == _T_807 ? 9'h36 : _GEN_95; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_98 = 8'h31 == _T_807 ? 1'h1 : _GEN_96; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_99 = 8'h31 == _T_807 ? 9'h65 : _GEN_97; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_100 = 8'h32 == _T_807 ? 1'h1 : _GEN_98; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_101 = 8'h32 == _T_807 ? 9'h69 : _GEN_99; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_102 = 8'h33 == _T_807 ? 1'h1 : _GEN_100; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_103 = 8'h33 == _T_807 ? 9'h6c : _GEN_101; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_104 = 8'h34 == _T_807 ? 1'h0 : _GEN_102; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_105 = 8'h34 == _T_807 ? 9'h0 : _GEN_103; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_106 = 8'h35 == _T_807 ? 1'h0 : _GEN_104; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_107 = 8'h35 == _T_807 ? 9'h0 : _GEN_105; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_108 = 8'h36 == _T_807 ? 1'h0 : _GEN_106; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_109 = 8'h36 == _T_807 ? 9'h0 : _GEN_107; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_110 = 8'h37 == _T_807 ? 1'h0 : _GEN_108; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_111 = 8'h37 == _T_807 ? 9'h0 : _GEN_109; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_112 = 8'h38 == _T_807 ? 1'h0 : _GEN_110; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_113 = 8'h38 == _T_807 ? 9'h0 : _GEN_111; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_114 = 8'h39 == _T_807 ? 1'h0 : _GEN_112; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_115 = 8'h39 == _T_807 ? 9'h0 : _GEN_113; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_116 = 8'h3a == _T_807 ? 1'h0 : _GEN_114; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_117 = 8'h3a == _T_807 ? 9'h0 : _GEN_115; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_118 = 8'h3b == _T_807 ? 1'h0 : _GEN_116; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_119 = 8'h3b == _T_807 ? 9'h0 : _GEN_117; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_120 = 8'h3c == _T_807 ? 1'h0 : _GEN_118; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_121 = 8'h3c == _T_807 ? 9'h0 : _GEN_119; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_122 = 8'h3d == _T_807 ? 1'h0 : _GEN_120; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_123 = 8'h3d == _T_807 ? 9'h0 : _GEN_121; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_124 = 8'h3e == _T_807 ? 1'h0 : _GEN_122; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_125 = 8'h3e == _T_807 ? 9'h0 : _GEN_123; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_126 = 8'h3f == _T_807 ? 1'h0 : _GEN_124; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_127 = 8'h3f == _T_807 ? 9'h0 : _GEN_125; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_128 = 8'h40 == _T_807 ? 1'h0 : _GEN_126; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_129 = 8'h40 == _T_807 ? 9'h0 : _GEN_127; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_130 = 8'h41 == _T_807 ? 1'h0 : _GEN_128; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_131 = 8'h41 == _T_807 ? 9'h0 : _GEN_129; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_132 = 8'h42 == _T_807 ? 1'h0 : _GEN_130; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_133 = 8'h42 == _T_807 ? 9'h0 : _GEN_131; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_134 = 8'h43 == _T_807 ? 1'h0 : _GEN_132; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_135 = 8'h43 == _T_807 ? 9'h0 : _GEN_133; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_136 = 8'h44 == _T_807 ? 1'h0 : _GEN_134; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_137 = 8'h44 == _T_807 ? 9'h0 : _GEN_135; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_138 = 8'h45 == _T_807 ? 1'h0 : _GEN_136; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_139 = 8'h45 == _T_807 ? 9'h0 : _GEN_137; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_140 = 8'h46 == _T_807 ? 1'h0 : _GEN_138; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_141 = 8'h46 == _T_807 ? 9'h0 : _GEN_139; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_142 = 8'h47 == _T_807 ? 1'h0 : _GEN_140; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_143 = 8'h47 == _T_807 ? 9'h0 : _GEN_141; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_144 = 8'h48 == _T_807 ? 1'h0 : _GEN_142; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_145 = 8'h48 == _T_807 ? 9'h0 : _GEN_143; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_146 = 8'h49 == _T_807 ? 1'h0 : _GEN_144; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_147 = 8'h49 == _T_807 ? 9'h0 : _GEN_145; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_148 = 8'h4a == _T_807 ? 1'h0 : _GEN_146; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_149 = 8'h4a == _T_807 ? 9'h0 : _GEN_147; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_150 = 8'h4b == _T_807 ? 1'h0 : _GEN_148; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_151 = 8'h4b == _T_807 ? 9'h0 : _GEN_149; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_152 = 8'h4c == _T_807 ? 1'h0 : _GEN_150; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_153 = 8'h4c == _T_807 ? 9'h0 : _GEN_151; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_154 = 8'h4d == _T_807 ? 1'h0 : _GEN_152; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_155 = 8'h4d == _T_807 ? 9'h0 : _GEN_153; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_156 = 8'h4e == _T_807 ? 1'h0 : _GEN_154; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_157 = 8'h4e == _T_807 ? 9'h0 : _GEN_155; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_158 = 8'h4f == _T_807 ? 1'h0 : _GEN_156; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_159 = 8'h4f == _T_807 ? 9'h0 : _GEN_157; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_160 = 8'h50 == _T_807 ? 1'h0 : _GEN_158; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_161 = 8'h50 == _T_807 ? 9'h0 : _GEN_159; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_162 = 8'h51 == _T_807 ? 1'h0 : _GEN_160; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_163 = 8'h51 == _T_807 ? 9'h0 : _GEN_161; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_164 = 8'h52 == _T_807 ? 1'h0 : _GEN_162; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_165 = 8'h52 == _T_807 ? 9'h0 : _GEN_163; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_166 = 8'h53 == _T_807 ? 1'h0 : _GEN_164; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_167 = 8'h53 == _T_807 ? 9'h0 : _GEN_165; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_168 = 8'h54 == _T_807 ? 1'h0 : _GEN_166; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_169 = 8'h54 == _T_807 ? 9'h0 : _GEN_167; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_170 = 8'h55 == _T_807 ? 1'h0 : _GEN_168; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_171 = 8'h55 == _T_807 ? 9'h0 : _GEN_169; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_172 = 8'h56 == _T_807 ? 1'h0 : _GEN_170; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_173 = 8'h56 == _T_807 ? 9'h0 : _GEN_171; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_174 = 8'h57 == _T_807 ? 1'h0 : _GEN_172; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_175 = 8'h57 == _T_807 ? 9'h0 : _GEN_173; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_176 = 8'h58 == _T_807 ? 1'h0 : _GEN_174; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_177 = 8'h58 == _T_807 ? 9'h0 : _GEN_175; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_178 = 8'h59 == _T_807 ? 1'h0 : _GEN_176; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_179 = 8'h59 == _T_807 ? 9'h0 : _GEN_177; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_180 = 8'h5a == _T_807 ? 1'h0 : _GEN_178; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_181 = 8'h5a == _T_807 ? 9'h0 : _GEN_179; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_182 = 8'h5b == _T_807 ? 1'h0 : _GEN_180; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_183 = 8'h5b == _T_807 ? 9'h0 : _GEN_181; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_184 = 8'h5c == _T_807 ? 1'h0 : _GEN_182; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_185 = 8'h5c == _T_807 ? 9'h0 : _GEN_183; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_186 = 8'h5d == _T_807 ? 1'h0 : _GEN_184; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_187 = 8'h5d == _T_807 ? 9'h0 : _GEN_185; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_188 = 8'h5e == _T_807 ? 1'h0 : _GEN_186; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_189 = 8'h5e == _T_807 ? 9'h0 : _GEN_187; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_190 = 8'h5f == _T_807 ? 1'h0 : _GEN_188; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_191 = 8'h5f == _T_807 ? 9'h0 : _GEN_189; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_192 = 8'h60 == _T_807 ? 1'h0 : _GEN_190; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_193 = 8'h60 == _T_807 ? 9'h0 : _GEN_191; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_194 = 8'h61 == _T_807 ? 1'h0 : _GEN_192; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_195 = 8'h61 == _T_807 ? 9'h0 : _GEN_193; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_196 = 8'h62 == _T_807 ? 1'h0 : _GEN_194; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_197 = 8'h62 == _T_807 ? 9'h0 : _GEN_195; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_198 = 8'h63 == _T_807 ? 1'h0 : _GEN_196; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_199 = 8'h63 == _T_807 ? 9'h0 : _GEN_197; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_200 = 8'h64 == _T_807 ? 1'h0 : _GEN_198; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_201 = 8'h64 == _T_807 ? 9'h0 : _GEN_199; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_202 = 8'h65 == _T_807 ? 1'h0 : _GEN_200; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_203 = 8'h65 == _T_807 ? 9'h0 : _GEN_201; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_204 = 8'h66 == _T_807 ? 1'h0 : _GEN_202; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_205 = 8'h66 == _T_807 ? 9'h0 : _GEN_203; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_206 = 8'h67 == _T_807 ? 1'h0 : _GEN_204; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_207 = 8'h67 == _T_807 ? 9'h0 : _GEN_205; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_208 = 8'h68 == _T_807 ? 1'h0 : _GEN_206; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_209 = 8'h68 == _T_807 ? 9'h0 : _GEN_207; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_210 = 8'h69 == _T_807 ? 1'h1 : _GEN_208; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_211 = 8'h69 == _T_807 ? 9'h30 : _GEN_209; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_212 = 8'h6a == _T_807 ? 1'h1 : _GEN_210; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_213 = 8'h6a == _T_807 ? 9'h32 : _GEN_211; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_214 = 8'h6b == _T_807 ? 1'h1 : _GEN_212; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_215 = 8'h6b == _T_807 ? 9'h35 : _GEN_213; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_216 = 8'h6c == _T_807 ? 1'h1 : _GEN_214; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_217 = 8'h6c == _T_807 ? 9'h61 : _GEN_215; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_218 = 8'h6d == _T_807 ? 1'h1 : _GEN_216; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_219 = 8'h6d == _T_807 ? 9'h66 : _GEN_217; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_220 = 8'h6e == _T_807 ? 1'h1 : _GEN_218; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_221 = 8'h6e == _T_807 ? 9'h6d : _GEN_219; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_222 = 8'h6f == _T_807 ? 1'h1 : _GEN_220; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_223 = 8'h6f == _T_807 ? 9'h6f : _GEN_221; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_224 = 8'h70 == _T_807 ? 1'h1 : _GEN_222; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_225 = 8'h70 == _T_807 ? 9'h72 : _GEN_223; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_226 = 8'h71 == _T_807 ? 1'h1 : _GEN_224; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_227 = 8'h71 == _T_807 ? 9'h73 : _GEN_225; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_228 = 8'h72 == _T_807 ? 1'h1 : _GEN_226; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_229 = 8'h72 == _T_807 ? 9'h78 : _GEN_227; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_230 = 8'h73 == _T_807 ? 1'h1 : _GEN_228; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_231 = 8'h73 == _T_807 ? 9'h101 : _GEN_229; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_232 = 8'h74 == _T_807 ? 1'h1 : _GEN_230; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_233 = 8'h74 == _T_807 ? 9'h102 : _GEN_231; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_234 = 8'h75 == _T_807 ? 1'h1 : _GEN_232; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_235 = 8'h75 == _T_807 ? 9'h116 : _GEN_233; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_236 = 8'h76 == _T_807 ? 1'h0 : _GEN_234; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_237 = 8'h76 == _T_807 ? 9'h0 : _GEN_235; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_238 = 8'h77 == _T_807 ? 1'h0 : _GEN_236; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_239 = 8'h77 == _T_807 ? 9'h0 : _GEN_237; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_240 = 8'h78 == _T_807 ? 1'h0 : _GEN_238; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_241 = 8'h78 == _T_807 ? 9'h0 : _GEN_239; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_242 = 8'h79 == _T_807 ? 1'h0 : _GEN_240; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_243 = 8'h79 == _T_807 ? 9'h0 : _GEN_241; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_244 = 8'h7a == _T_807 ? 1'h0 : _GEN_242; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_245 = 8'h7a == _T_807 ? 9'h0 : _GEN_243; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_246 = 8'h7b == _T_807 ? 1'h0 : _GEN_244; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_247 = 8'h7b == _T_807 ? 9'h0 : _GEN_245; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_248 = 8'h7c == _T_807 ? 1'h0 : _GEN_246; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_249 = 8'h7c == _T_807 ? 9'h0 : _GEN_247; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_250 = 8'h7d == _T_807 ? 1'h0 : _GEN_248; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_251 = 8'h7d == _T_807 ? 9'h0 : _GEN_249; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_252 = 8'h7e == _T_807 ? 1'h0 : _GEN_250; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_253 = 8'h7e == _T_807 ? 9'h0 : _GEN_251; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_254 = 8'h7f == _T_807 ? 1'h0 : _GEN_252; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_255 = 8'h7f == _T_807 ? 9'h0 : _GEN_253; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_256 = 8'h80 == _T_807 ? 1'h0 : _GEN_254; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_257 = 8'h80 == _T_807 ? 9'h0 : _GEN_255; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_258 = 8'h81 == _T_807 ? 1'h0 : _GEN_256; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_259 = 8'h81 == _T_807 ? 9'h0 : _GEN_257; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_260 = 8'h82 == _T_807 ? 1'h0 : _GEN_258; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_261 = 8'h82 == _T_807 ? 9'h0 : _GEN_259; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_262 = 8'h83 == _T_807 ? 1'h0 : _GEN_260; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_263 = 8'h83 == _T_807 ? 9'h0 : _GEN_261; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_264 = 8'h84 == _T_807 ? 1'h0 : _GEN_262; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_265 = 8'h84 == _T_807 ? 9'h0 : _GEN_263; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_266 = 8'h85 == _T_807 ? 1'h0 : _GEN_264; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_267 = 8'h85 == _T_807 ? 9'h0 : _GEN_265; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_268 = 8'h86 == _T_807 ? 1'h0 : _GEN_266; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_269 = 8'h86 == _T_807 ? 9'h0 : _GEN_267; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_270 = 8'h87 == _T_807 ? 1'h0 : _GEN_268; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_271 = 8'h87 == _T_807 ? 9'h0 : _GEN_269; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_272 = 8'h88 == _T_807 ? 1'h0 : _GEN_270; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_273 = 8'h88 == _T_807 ? 9'h0 : _GEN_271; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_274 = 8'h89 == _T_807 ? 1'h0 : _GEN_272; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_275 = 8'h89 == _T_807 ? 9'h0 : _GEN_273; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_276 = 8'h8a == _T_807 ? 1'h0 : _GEN_274; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_277 = 8'h8a == _T_807 ? 9'h0 : _GEN_275; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_278 = 8'h8b == _T_807 ? 1'h0 : _GEN_276; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_279 = 8'h8b == _T_807 ? 9'h0 : _GEN_277; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_280 = 8'h8c == _T_807 ? 1'h0 : _GEN_278; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_281 = 8'h8c == _T_807 ? 9'h0 : _GEN_279; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_282 = 8'h8d == _T_807 ? 1'h0 : _GEN_280; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_283 = 8'h8d == _T_807 ? 9'h0 : _GEN_281; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_284 = 8'h8e == _T_807 ? 1'h0 : _GEN_282; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_285 = 8'h8e == _T_807 ? 9'h0 : _GEN_283; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_286 = 8'h8f == _T_807 ? 1'h0 : _GEN_284; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_287 = 8'h8f == _T_807 ? 9'h0 : _GEN_285; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_288 = 8'h90 == _T_807 ? 1'h0 : _GEN_286; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_289 = 8'h90 == _T_807 ? 9'h0 : _GEN_287; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_290 = 8'h91 == _T_807 ? 1'h0 : _GEN_288; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_291 = 8'h91 == _T_807 ? 9'h0 : _GEN_289; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_292 = 8'h92 == _T_807 ? 1'h0 : _GEN_290; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_293 = 8'h92 == _T_807 ? 9'h0 : _GEN_291; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_294 = 8'h93 == _T_807 ? 1'h0 : _GEN_292; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_295 = 8'h93 == _T_807 ? 9'h0 : _GEN_293; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_296 = 8'h94 == _T_807 ? 1'h0 : _GEN_294; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_297 = 8'h94 == _T_807 ? 9'h0 : _GEN_295; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_298 = 8'h95 == _T_807 ? 1'h0 : _GEN_296; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_299 = 8'h95 == _T_807 ? 9'h0 : _GEN_297; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_300 = 8'h96 == _T_807 ? 1'h0 : _GEN_298; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_301 = 8'h96 == _T_807 ? 9'h0 : _GEN_299; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_302 = 8'h97 == _T_807 ? 1'h0 : _GEN_300; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_303 = 8'h97 == _T_807 ? 9'h0 : _GEN_301; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_304 = 8'h98 == _T_807 ? 1'h0 : _GEN_302; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_305 = 8'h98 == _T_807 ? 9'h0 : _GEN_303; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_306 = 8'h99 == _T_807 ? 1'h0 : _GEN_304; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_307 = 8'h99 == _T_807 ? 9'h0 : _GEN_305; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_308 = 8'h9a == _T_807 ? 1'h0 : _GEN_306; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_309 = 8'h9a == _T_807 ? 9'h0 : _GEN_307; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_310 = 8'h9b == _T_807 ? 1'h0 : _GEN_308; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_311 = 8'h9b == _T_807 ? 9'h0 : _GEN_309; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_312 = 8'h9c == _T_807 ? 1'h0 : _GEN_310; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_313 = 8'h9c == _T_807 ? 9'h0 : _GEN_311; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_314 = 8'h9d == _T_807 ? 1'h0 : _GEN_312; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_315 = 8'h9d == _T_807 ? 9'h0 : _GEN_313; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_316 = 8'h9e == _T_807 ? 1'h0 : _GEN_314; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_317 = 8'h9e == _T_807 ? 9'h0 : _GEN_315; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_318 = 8'h9f == _T_807 ? 1'h0 : _GEN_316; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_319 = 8'h9f == _T_807 ? 9'h0 : _GEN_317; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_320 = 8'ha0 == _T_807 ? 1'h0 : _GEN_318; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_321 = 8'ha0 == _T_807 ? 9'h0 : _GEN_319; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_322 = 8'ha1 == _T_807 ? 1'h0 : _GEN_320; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_323 = 8'ha1 == _T_807 ? 9'h0 : _GEN_321; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_324 = 8'ha2 == _T_807 ? 1'h0 : _GEN_322; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_325 = 8'ha2 == _T_807 ? 9'h0 : _GEN_323; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_326 = 8'ha3 == _T_807 ? 1'h0 : _GEN_324; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_327 = 8'ha3 == _T_807 ? 9'h0 : _GEN_325; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_328 = 8'ha4 == _T_807 ? 1'h0 : _GEN_326; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_329 = 8'ha4 == _T_807 ? 9'h0 : _GEN_327; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_330 = 8'ha5 == _T_807 ? 1'h0 : _GEN_328; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_331 = 8'ha5 == _T_807 ? 9'h0 : _GEN_329; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_332 = 8'ha6 == _T_807 ? 1'h0 : _GEN_330; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_333 = 8'ha6 == _T_807 ? 9'h0 : _GEN_331; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_334 = 8'ha7 == _T_807 ? 1'h0 : _GEN_332; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_335 = 8'ha7 == _T_807 ? 9'h0 : _GEN_333; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_336 = 8'ha8 == _T_807 ? 1'h0 : _GEN_334; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_337 = 8'ha8 == _T_807 ? 9'h0 : _GEN_335; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_338 = 8'ha9 == _T_807 ? 1'h0 : _GEN_336; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_339 = 8'ha9 == _T_807 ? 9'h0 : _GEN_337; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_340 = 8'haa == _T_807 ? 1'h0 : _GEN_338; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_341 = 8'haa == _T_807 ? 9'h0 : _GEN_339; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_342 = 8'hab == _T_807 ? 1'h0 : _GEN_340; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_343 = 8'hab == _T_807 ? 9'h0 : _GEN_341; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_344 = 8'hac == _T_807 ? 1'h0 : _GEN_342; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_345 = 8'hac == _T_807 ? 9'h0 : _GEN_343; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_346 = 8'had == _T_807 ? 1'h0 : _GEN_344; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_347 = 8'had == _T_807 ? 9'h0 : _GEN_345; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_348 = 8'hae == _T_807 ? 1'h0 : _GEN_346; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_349 = 8'hae == _T_807 ? 9'h0 : _GEN_347; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_350 = 8'haf == _T_807 ? 1'h0 : _GEN_348; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_351 = 8'haf == _T_807 ? 9'h0 : _GEN_349; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_352 = 8'hb0 == _T_807 ? 1'h0 : _GEN_350; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_353 = 8'hb0 == _T_807 ? 9'h0 : _GEN_351; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_354 = 8'hb1 == _T_807 ? 1'h0 : _GEN_352; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_355 = 8'hb1 == _T_807 ? 9'h0 : _GEN_353; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_356 = 8'hb2 == _T_807 ? 1'h0 : _GEN_354; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_357 = 8'hb2 == _T_807 ? 9'h0 : _GEN_355; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_358 = 8'hb3 == _T_807 ? 1'h0 : _GEN_356; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_359 = 8'hb3 == _T_807 ? 9'h0 : _GEN_357; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_360 = 8'hb4 == _T_807 ? 1'h0 : _GEN_358; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_361 = 8'hb4 == _T_807 ? 9'h0 : _GEN_359; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_362 = 8'hb5 == _T_807 ? 1'h0 : _GEN_360; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_363 = 8'hb5 == _T_807 ? 9'h0 : _GEN_361; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_364 = 8'hb6 == _T_807 ? 1'h0 : _GEN_362; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_365 = 8'hb6 == _T_807 ? 9'h0 : _GEN_363; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_366 = 8'hb7 == _T_807 ? 1'h0 : _GEN_364; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_367 = 8'hb7 == _T_807 ? 9'h0 : _GEN_365; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_368 = 8'hb8 == _T_807 ? 1'h0 : _GEN_366; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_369 = 8'hb8 == _T_807 ? 9'h0 : _GEN_367; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_370 = 8'hb9 == _T_807 ? 1'h0 : _GEN_368; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_371 = 8'hb9 == _T_807 ? 9'h0 : _GEN_369; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_372 = 8'hba == _T_807 ? 1'h0 : _GEN_370; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_373 = 8'hba == _T_807 ? 9'h0 : _GEN_371; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_374 = 8'hbb == _T_807 ? 1'h0 : _GEN_372; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_375 = 8'hbb == _T_807 ? 9'h0 : _GEN_373; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_376 = 8'hbc == _T_807 ? 1'h0 : _GEN_374; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_377 = 8'hbc == _T_807 ? 9'h0 : _GEN_375; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_378 = 8'hbd == _T_807 ? 1'h0 : _GEN_376; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_379 = 8'hbd == _T_807 ? 9'h0 : _GEN_377; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_380 = 8'hbe == _T_807 ? 1'h0 : _GEN_378; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_381 = 8'hbe == _T_807 ? 9'h0 : _GEN_379; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_382 = 8'hbf == _T_807 ? 1'h0 : _GEN_380; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_383 = 8'hbf == _T_807 ? 9'h0 : _GEN_381; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_384 = 8'hc0 == _T_807 ? 1'h0 : _GEN_382; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_385 = 8'hc0 == _T_807 ? 9'h0 : _GEN_383; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_386 = 8'hc1 == _T_807 ? 1'h0 : _GEN_384; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_387 = 8'hc1 == _T_807 ? 9'h0 : _GEN_385; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_388 = 8'hc2 == _T_807 ? 1'h0 : _GEN_386; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_389 = 8'hc2 == _T_807 ? 9'h0 : _GEN_387; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_390 = 8'hc3 == _T_807 ? 1'h0 : _GEN_388; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_391 = 8'hc3 == _T_807 ? 9'h0 : _GEN_389; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_392 = 8'hc4 == _T_807 ? 1'h0 : _GEN_390; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_393 = 8'hc4 == _T_807 ? 9'h0 : _GEN_391; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_394 = 8'hc5 == _T_807 ? 1'h0 : _GEN_392; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_395 = 8'hc5 == _T_807 ? 9'h0 : _GEN_393; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_396 = 8'hc6 == _T_807 ? 1'h0 : _GEN_394; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_397 = 8'hc6 == _T_807 ? 9'h0 : _GEN_395; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_398 = 8'hc7 == _T_807 ? 1'h0 : _GEN_396; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_399 = 8'hc7 == _T_807 ? 9'h0 : _GEN_397; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_400 = 8'hc8 == _T_807 ? 1'h0 : _GEN_398; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_401 = 8'hc8 == _T_807 ? 9'h0 : _GEN_399; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_402 = 8'hc9 == _T_807 ? 1'h0 : _GEN_400; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_403 = 8'hc9 == _T_807 ? 9'h0 : _GEN_401; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_404 = 8'hca == _T_807 ? 1'h0 : _GEN_402; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_405 = 8'hca == _T_807 ? 9'h0 : _GEN_403; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_406 = 8'hcb == _T_807 ? 1'h0 : _GEN_404; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_407 = 8'hcb == _T_807 ? 9'h0 : _GEN_405; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_408 = 8'hcc == _T_807 ? 1'h0 : _GEN_406; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_409 = 8'hcc == _T_807 ? 9'h0 : _GEN_407; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_410 = 8'hcd == _T_807 ? 1'h0 : _GEN_408; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_411 = 8'hcd == _T_807 ? 9'h0 : _GEN_409; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_412 = 8'hce == _T_807 ? 1'h0 : _GEN_410; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_413 = 8'hce == _T_807 ? 9'h0 : _GEN_411; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_414 = 8'hcf == _T_807 ? 1'h0 : _GEN_412; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_415 = 8'hcf == _T_807 ? 9'h0 : _GEN_413; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_416 = 8'hd0 == _T_807 ? 1'h0 : _GEN_414; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_417 = 8'hd0 == _T_807 ? 9'h0 : _GEN_415; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_418 = 8'hd1 == _T_807 ? 1'h0 : _GEN_416; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_419 = 8'hd1 == _T_807 ? 9'h0 : _GEN_417; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_420 = 8'hd2 == _T_807 ? 1'h0 : _GEN_418; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_421 = 8'hd2 == _T_807 ? 9'h0 : _GEN_419; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_422 = 8'hd3 == _T_807 ? 1'h0 : _GEN_420; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_423 = 8'hd3 == _T_807 ? 9'h0 : _GEN_421; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_424 = 8'hd4 == _T_807 ? 1'h0 : _GEN_422; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_425 = 8'hd4 == _T_807 ? 9'h0 : _GEN_423; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_426 = 8'hd5 == _T_807 ? 1'h0 : _GEN_424; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_427 = 8'hd5 == _T_807 ? 9'h0 : _GEN_425; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_428 = 8'hd6 == _T_807 ? 1'h0 : _GEN_426; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_429 = 8'hd6 == _T_807 ? 9'h0 : _GEN_427; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_430 = 8'hd7 == _T_807 ? 1'h0 : _GEN_428; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_431 = 8'hd7 == _T_807 ? 9'h0 : _GEN_429; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_432 = 8'hd8 == _T_807 ? 1'h0 : _GEN_430; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_433 = 8'hd8 == _T_807 ? 9'h0 : _GEN_431; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_434 = 8'hd9 == _T_807 ? 1'h0 : _GEN_432; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_435 = 8'hd9 == _T_807 ? 9'h0 : _GEN_433; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_436 = 8'hda == _T_807 ? 1'h0 : _GEN_434; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_437 = 8'hda == _T_807 ? 9'h0 : _GEN_435; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_438 = 8'hdb == _T_807 ? 1'h0 : _GEN_436; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_439 = 8'hdb == _T_807 ? 9'h0 : _GEN_437; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_440 = 8'hdc == _T_807 ? 1'h0 : _GEN_438; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_441 = 8'hdc == _T_807 ? 9'h0 : _GEN_439; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_442 = 8'hdd == _T_807 ? 1'h0 : _GEN_440; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_443 = 8'hdd == _T_807 ? 9'h0 : _GEN_441; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_444 = 8'hde == _T_807 ? 1'h0 : _GEN_442; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_445 = 8'hde == _T_807 ? 9'h0 : _GEN_443; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_446 = 8'hdf == _T_807 ? 1'h0 : _GEN_444; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_447 = 8'hdf == _T_807 ? 9'h0 : _GEN_445; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_448 = 8'he0 == _T_807 ? 1'h0 : _GEN_446; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_449 = 8'he0 == _T_807 ? 9'h0 : _GEN_447; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_450 = 8'he1 == _T_807 ? 1'h0 : _GEN_448; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_451 = 8'he1 == _T_807 ? 9'h0 : _GEN_449; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_452 = 8'he2 == _T_807 ? 1'h0 : _GEN_450; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_453 = 8'he2 == _T_807 ? 9'h0 : _GEN_451; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_454 = 8'he3 == _T_807 ? 1'h0 : _GEN_452; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_455 = 8'he3 == _T_807 ? 9'h0 : _GEN_453; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_456 = 8'he4 == _T_807 ? 1'h0 : _GEN_454; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_457 = 8'he4 == _T_807 ? 9'h0 : _GEN_455; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_458 = 8'he5 == _T_807 ? 1'h0 : _GEN_456; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_459 = 8'he5 == _T_807 ? 9'h0 : _GEN_457; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_460 = 8'he6 == _T_807 ? 1'h0 : _GEN_458; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_461 = 8'he6 == _T_807 ? 9'h0 : _GEN_459; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_462 = 8'he7 == _T_807 ? 1'h0 : _GEN_460; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_463 = 8'he7 == _T_807 ? 9'h0 : _GEN_461; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_464 = 8'he8 == _T_807 ? 1'h0 : _GEN_462; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_465 = 8'he8 == _T_807 ? 9'h0 : _GEN_463; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_466 = 8'he9 == _T_807 ? 1'h0 : _GEN_464; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_467 = 8'he9 == _T_807 ? 9'h0 : _GEN_465; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_468 = 8'hea == _T_807 ? 1'h0 : _GEN_466; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_469 = 8'hea == _T_807 ? 9'h0 : _GEN_467; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_470 = 8'heb == _T_807 ? 1'h0 : _GEN_468; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_471 = 8'heb == _T_807 ? 9'h0 : _GEN_469; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_472 = 8'hec == _T_807 ? 1'h0 : _GEN_470; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_473 = 8'hec == _T_807 ? 9'h0 : _GEN_471; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_474 = 8'hed == _T_807 ? 1'h1 : _GEN_472; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_475 = 8'hed == _T_807 ? 9'h21 : _GEN_473; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_476 = 8'hee == _T_807 ? 1'h1 : _GEN_474; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_477 = 8'hee == _T_807 ? 9'h2e : _GEN_475; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_478 = 8'hef == _T_807 ? 1'h1 : _GEN_476; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_479 = 8'hef == _T_807 ? 9'h37 : _GEN_477; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_480 = 8'hf0 == _T_807 ? 1'h1 : _GEN_478; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_481 = 8'hf0 == _T_807 ? 9'h48 : _GEN_479; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_482 = 8'hf1 == _T_807 ? 1'h1 : _GEN_480; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_483 = 8'hf1 == _T_807 ? 9'h67 : _GEN_481; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_484 = 8'hf2 == _T_807 ? 1'h1 : _GEN_482; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_485 = 8'hf2 == _T_807 ? 9'h6a : _GEN_483; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_486 = 8'hf3 == _T_807 ? 1'h1 : _GEN_484; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_487 = 8'hf3 == _T_807 ? 9'h6e : _GEN_485; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_488 = 8'hf4 == _T_807 ? 1'h1 : _GEN_486; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_489 = 8'hf4 == _T_807 ? 9'h70 : _GEN_487; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_490 = 8'hf5 == _T_807 ? 1'h1 : _GEN_488; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_491 = 8'hf5 == _T_807 ? 9'h75 : _GEN_489; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_492 = 8'hf6 == _T_807 ? 1'h1 : _GEN_490; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_493 = 8'hf6 == _T_807 ? 9'h100 : _GEN_491; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_494 = 8'hf7 == _T_807 ? 1'h1 : _GEN_492; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_495 = 8'hf7 == _T_807 ? 9'h104 : _GEN_493; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_496 = 8'hf8 == _T_807 ? 1'h1 : _GEN_494; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_497 = 8'hf8 == _T_807 ? 9'h106 : _GEN_495; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_498 = 8'hf9 == _T_807 ? 1'h1 : _GEN_496; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_499 = 8'hf9 == _T_807 ? 9'h108 : _GEN_497; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_500 = 8'hfa == _T_807 ? 1'h1 : _GEN_498; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_501 = 8'hfa == _T_807 ? 9'h109 : _GEN_499; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_502 = 8'hfb == _T_807 ? 1'h1 : _GEN_500; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_503 = 8'hfb == _T_807 ? 9'h10f : _GEN_501; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_504 = 8'hfc == _T_807 ? 1'h1 : _GEN_502; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_505 = 8'hfc == _T_807 ? 9'h110 : _GEN_503; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_506 = 8'hfd == _T_807 ? 1'h1 : _GEN_504; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_507 = 8'hfd == _T_807 ? 9'h118 : _GEN_505; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_508 = 8'hfe == _T_807 ? 1'h1 : _GEN_506; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_509 = 8'hfe == _T_807 ? 9'h11a : _GEN_507; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_1530 = _GEN_508 ? 11'h0 : _T_805; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_1531 = _GEN_508 ? 1'h0 : 1'h1; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_1532 = _GEN_508 ? _GEN_509 : data_reg; // @[GunzipHuffDecoder.scala 60:43:@564.10]
  assign _GEN_1535 = io_enable ? _GEN_1531 : 1'h0; // @[GunzipHuffDecoder.scala 55:29:@555.8]
  assign _GEN_1536 = io_enable ? _GEN_1530 : 11'h0; // @[GunzipHuffDecoder.scala 55:29:@555.8]
  assign _GEN_1537 = io_enable ? _GEN_1532 : data_reg; // @[GunzipHuffDecoder.scala 55:29:@555.8]
  assign _GEN_1539 = io_enable ? _GEN_508 : 1'h0; // @[GunzipHuffDecoder.scala 55:29:@555.8]
  assign _GEN_1540 = _T_794 ? 1'h0 : _GEN_1535; // @[GunzipHuffDecoder.scala 52:46:@547.6]
  assign _GEN_1541 = _T_794 ? {{2'd0}, lit_idx} : _GEN_1536; // @[GunzipHuffDecoder.scala 52:46:@547.6]
  assign _GEN_1542 = _T_794 ? data_reg : _GEN_1537; // @[GunzipHuffDecoder.scala 52:46:@547.6]
  assign _GEN_1544 = _T_794 ? 1'h0 : _GEN_1539; // @[GunzipHuffDecoder.scala 52:46:@547.6]
  assign _GEN_1546 = io_data_in_valid ? _GEN_1541 : {{2'd0}, lit_idx}; // @[GunzipHuffDecoder.scala 51:27:@545.4]
  assign io_data_in_ready = io_data_in_valid ? _GEN_1540 : 1'h0; // @[GunzipHuffDecoder.scala 46:20:@542.4 GunzipHuffDecoder.scala 56:24:@556.10 GunzipHuffDecoder.scala 62:26:@566.12]
  assign io_data = io_data_in_valid ? _GEN_1542 : data_reg; // @[GunzipHuffDecoder.scala 48:11:@543.4 GunzipHuffDecoder.scala 63:17:@568.12]
  assign io_valid = io_data_in_valid ? _GEN_1544 : 1'h0; // @[GunzipHuffDecoder.scala 49:12:@544.4 GunzipHuffDecoder.scala 65:18:@571.12]
  assign _GEN_1551 = io_data_in_valid & _T_794; // @[GunzipHuffDecoder.scala 54:13:@551.10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lit_idx = _RAND_0[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  data_reg = _RAND_1[8:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      lit_idx <= 9'h0;
    end else begin
      lit_idx <= _GEN_1546[8:0];
    end
    if (io_data_in_valid) begin
      if (!(_T_794)) begin
        if (io_enable) begin
          if (_GEN_508) begin
            if (8'hfe == _T_807) begin
              data_reg <= 9'h11a;
            end else begin
              if (8'hfd == _T_807) begin
                data_reg <= 9'h118;
              end else begin
                if (8'hfc == _T_807) begin
                  data_reg <= 9'h110;
                end else begin
                  if (8'hfb == _T_807) begin
                    data_reg <= 9'h10f;
                  end else begin
                    if (8'hfa == _T_807) begin
                      data_reg <= 9'h109;
                    end else begin
                      if (8'hf9 == _T_807) begin
                        data_reg <= 9'h108;
                      end else begin
                        if (8'hf8 == _T_807) begin
                          data_reg <= 9'h106;
                        end else begin
                          if (8'hf7 == _T_807) begin
                            data_reg <= 9'h104;
                          end else begin
                            if (8'hf6 == _T_807) begin
                              data_reg <= 9'h100;
                            end else begin
                              if (8'hf5 == _T_807) begin
                                data_reg <= 9'h75;
                              end else begin
                                if (8'hf4 == _T_807) begin
                                  data_reg <= 9'h70;
                                end else begin
                                  if (8'hf3 == _T_807) begin
                                    data_reg <= 9'h6e;
                                  end else begin
                                    if (8'hf2 == _T_807) begin
                                      data_reg <= 9'h6a;
                                    end else begin
                                      if (8'hf1 == _T_807) begin
                                        data_reg <= 9'h67;
                                      end else begin
                                        if (8'hf0 == _T_807) begin
                                          data_reg <= 9'h48;
                                        end else begin
                                          if (8'hef == _T_807) begin
                                            data_reg <= 9'h37;
                                          end else begin
                                            if (8'hee == _T_807) begin
                                              data_reg <= 9'h2e;
                                            end else begin
                                              if (8'hed == _T_807) begin
                                                data_reg <= 9'h21;
                                              end else begin
                                                if (8'hec == _T_807) begin
                                                  data_reg <= 9'h0;
                                                end else begin
                                                  if (8'heb == _T_807) begin
                                                    data_reg <= 9'h0;
                                                  end else begin
                                                    if (8'hea == _T_807) begin
                                                      data_reg <= 9'h0;
                                                    end else begin
                                                      if (8'he9 == _T_807) begin
                                                        data_reg <= 9'h0;
                                                      end else begin
                                                        if (8'he8 == _T_807) begin
                                                          data_reg <= 9'h0;
                                                        end else begin
                                                          if (8'he7 == _T_807) begin
                                                            data_reg <= 9'h0;
                                                          end else begin
                                                            if (8'he6 == _T_807) begin
                                                              data_reg <= 9'h0;
                                                            end else begin
                                                              if (8'he5 == _T_807) begin
                                                                data_reg <= 9'h0;
                                                              end else begin
                                                                if (8'he4 == _T_807) begin
                                                                  data_reg <= 9'h0;
                                                                end else begin
                                                                  if (8'he3 == _T_807) begin
                                                                    data_reg <= 9'h0;
                                                                  end else begin
                                                                    if (8'he2 == _T_807) begin
                                                                      data_reg <= 9'h0;
                                                                    end else begin
                                                                      if (8'he1 == _T_807) begin
                                                                        data_reg <= 9'h0;
                                                                      end else begin
                                                                        if (8'he0 == _T_807) begin
                                                                          data_reg <= 9'h0;
                                                                        end else begin
                                                                          if (8'hdf == _T_807) begin
                                                                            data_reg <= 9'h0;
                                                                          end else begin
                                                                            if (8'hde == _T_807) begin
                                                                              data_reg <= 9'h0;
                                                                            end else begin
                                                                              if (8'hdd == _T_807) begin
                                                                                data_reg <= 9'h0;
                                                                              end else begin
                                                                                if (8'hdc == _T_807) begin
                                                                                  data_reg <= 9'h0;
                                                                                end else begin
                                                                                  if (8'hdb == _T_807) begin
                                                                                    data_reg <= 9'h0;
                                                                                  end else begin
                                                                                    if (8'hda == _T_807) begin
                                                                                      data_reg <= 9'h0;
                                                                                    end else begin
                                                                                      if (8'hd9 == _T_807) begin
                                                                                        data_reg <= 9'h0;
                                                                                      end else begin
                                                                                        if (8'hd8 == _T_807) begin
                                                                                          data_reg <= 9'h0;
                                                                                        end else begin
                                                                                          if (8'hd7 == _T_807) begin
                                                                                            data_reg <= 9'h0;
                                                                                          end else begin
                                                                                            if (8'hd6 == _T_807) begin
                                                                                              data_reg <= 9'h0;
                                                                                            end else begin
                                                                                              if (8'hd5 == _T_807) begin
                                                                                                data_reg <= 9'h0;
                                                                                              end else begin
                                                                                                if (8'hd4 == _T_807) begin
                                                                                                  data_reg <= 9'h0;
                                                                                                end else begin
                                                                                                  if (8'hd3 == _T_807) begin
                                                                                                    data_reg <= 9'h0;
                                                                                                  end else begin
                                                                                                    if (8'hd2 == _T_807) begin
                                                                                                      data_reg <= 9'h0;
                                                                                                    end else begin
                                                                                                      if (8'hd1 == _T_807) begin
                                                                                                        data_reg <= 9'h0;
                                                                                                      end else begin
                                                                                                        if (8'hd0 == _T_807) begin
                                                                                                          data_reg <= 9'h0;
                                                                                                        end else begin
                                                                                                          if (8'hcf == _T_807) begin
                                                                                                            data_reg <= 9'h0;
                                                                                                          end else begin
                                                                                                            if (8'hce == _T_807) begin
                                                                                                              data_reg <= 9'h0;
                                                                                                            end else begin
                                                                                                              if (8'hcd == _T_807) begin
                                                                                                                data_reg <= 9'h0;
                                                                                                              end else begin
                                                                                                                if (8'hcc == _T_807) begin
                                                                                                                  data_reg <= 9'h0;
                                                                                                                end else begin
                                                                                                                  if (8'hcb == _T_807) begin
                                                                                                                    data_reg <= 9'h0;
                                                                                                                  end else begin
                                                                                                                    if (8'hca == _T_807) begin
                                                                                                                      data_reg <= 9'h0;
                                                                                                                    end else begin
                                                                                                                      if (8'hc9 == _T_807) begin
                                                                                                                        data_reg <= 9'h0;
                                                                                                                      end else begin
                                                                                                                        if (8'hc8 == _T_807) begin
                                                                                                                          data_reg <= 9'h0;
                                                                                                                        end else begin
                                                                                                                          if (8'hc7 == _T_807) begin
                                                                                                                            data_reg <= 9'h0;
                                                                                                                          end else begin
                                                                                                                            if (8'hc6 == _T_807) begin
                                                                                                                              data_reg <= 9'h0;
                                                                                                                            end else begin
                                                                                                                              if (8'hc5 == _T_807) begin
                                                                                                                                data_reg <= 9'h0;
                                                                                                                              end else begin
                                                                                                                                if (8'hc4 == _T_807) begin
                                                                                                                                  data_reg <= 9'h0;
                                                                                                                                end else begin
                                                                                                                                  if (8'hc3 == _T_807) begin
                                                                                                                                    data_reg <= 9'h0;
                                                                                                                                  end else begin
                                                                                                                                    if (8'hc2 == _T_807) begin
                                                                                                                                      data_reg <= 9'h0;
                                                                                                                                    end else begin
                                                                                                                                      if (8'hc1 == _T_807) begin
                                                                                                                                        data_reg <= 9'h0;
                                                                                                                                      end else begin
                                                                                                                                        if (8'hc0 == _T_807) begin
                                                                                                                                          data_reg <= 9'h0;
                                                                                                                                        end else begin
                                                                                                                                          if (8'hbf == _T_807) begin
                                                                                                                                            data_reg <= 9'h0;
                                                                                                                                          end else begin
                                                                                                                                            if (8'hbe == _T_807) begin
                                                                                                                                              data_reg <= 9'h0;
                                                                                                                                            end else begin
                                                                                                                                              if (8'hbd == _T_807) begin
                                                                                                                                                data_reg <= 9'h0;
                                                                                                                                              end else begin
                                                                                                                                                if (8'hbc == _T_807) begin
                                                                                                                                                  data_reg <= 9'h0;
                                                                                                                                                end else begin
                                                                                                                                                  if (8'hbb == _T_807) begin
                                                                                                                                                    data_reg <= 9'h0;
                                                                                                                                                  end else begin
                                                                                                                                                    if (8'hba == _T_807) begin
                                                                                                                                                      data_reg <= 9'h0;
                                                                                                                                                    end else begin
                                                                                                                                                      if (8'hb9 == _T_807) begin
                                                                                                                                                        data_reg <= 9'h0;
                                                                                                                                                      end else begin
                                                                                                                                                        if (8'hb8 == _T_807) begin
                                                                                                                                                          data_reg <= 9'h0;
                                                                                                                                                        end else begin
                                                                                                                                                          if (8'hb7 == _T_807) begin
                                                                                                                                                            data_reg <= 9'h0;
                                                                                                                                                          end else begin
                                                                                                                                                            if (8'hb6 == _T_807) begin
                                                                                                                                                              data_reg <= 9'h0;
                                                                                                                                                            end else begin
                                                                                                                                                              if (8'hb5 == _T_807) begin
                                                                                                                                                                data_reg <= 9'h0;
                                                                                                                                                              end else begin
                                                                                                                                                                if (8'hb4 == _T_807) begin
                                                                                                                                                                  data_reg <= 9'h0;
                                                                                                                                                                end else begin
                                                                                                                                                                  if (8'hb3 == _T_807) begin
                                                                                                                                                                    data_reg <= 9'h0;
                                                                                                                                                                  end else begin
                                                                                                                                                                    if (8'hb2 == _T_807) begin
                                                                                                                                                                      data_reg <= 9'h0;
                                                                                                                                                                    end else begin
                                                                                                                                                                      if (8'hb1 == _T_807) begin
                                                                                                                                                                        data_reg <= 9'h0;
                                                                                                                                                                      end else begin
                                                                                                                                                                        if (8'hb0 == _T_807) begin
                                                                                                                                                                          data_reg <= 9'h0;
                                                                                                                                                                        end else begin
                                                                                                                                                                          if (8'haf == _T_807) begin
                                                                                                                                                                            data_reg <= 9'h0;
                                                                                                                                                                          end else begin
                                                                                                                                                                            if (8'hae == _T_807) begin
                                                                                                                                                                              data_reg <= 9'h0;
                                                                                                                                                                            end else begin
                                                                                                                                                                              if (8'had == _T_807) begin
                                                                                                                                                                                data_reg <= 9'h0;
                                                                                                                                                                              end else begin
                                                                                                                                                                                if (8'hac == _T_807) begin
                                                                                                                                                                                  data_reg <= 9'h0;
                                                                                                                                                                                end else begin
                                                                                                                                                                                  if (8'hab == _T_807) begin
                                                                                                                                                                                    data_reg <= 9'h0;
                                                                                                                                                                                  end else begin
                                                                                                                                                                                    if (8'haa == _T_807) begin
                                                                                                                                                                                      data_reg <= 9'h0;
                                                                                                                                                                                    end else begin
                                                                                                                                                                                      if (8'ha9 == _T_807) begin
                                                                                                                                                                                        data_reg <= 9'h0;
                                                                                                                                                                                      end else begin
                                                                                                                                                                                        if (8'ha8 == _T_807) begin
                                                                                                                                                                                          data_reg <= 9'h0;
                                                                                                                                                                                        end else begin
                                                                                                                                                                                          if (8'ha7 == _T_807) begin
                                                                                                                                                                                            data_reg <= 9'h0;
                                                                                                                                                                                          end else begin
                                                                                                                                                                                            if (8'ha6 == _T_807) begin
                                                                                                                                                                                              data_reg <= 9'h0;
                                                                                                                                                                                            end else begin
                                                                                                                                                                                              if (8'ha5 == _T_807) begin
                                                                                                                                                                                                data_reg <= 9'h0;
                                                                                                                                                                                              end else begin
                                                                                                                                                                                                if (8'ha4 == _T_807) begin
                                                                                                                                                                                                  data_reg <= 9'h0;
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                  if (8'ha3 == _T_807) begin
                                                                                                                                                                                                    data_reg <= 9'h0;
                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                    if (8'ha2 == _T_807) begin
                                                                                                                                                                                                      data_reg <= 9'h0;
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                      if (8'ha1 == _T_807) begin
                                                                                                                                                                                                        data_reg <= 9'h0;
                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                        if (8'ha0 == _T_807) begin
                                                                                                                                                                                                          data_reg <= 9'h0;
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                          if (8'h9f == _T_807) begin
                                                                                                                                                                                                            data_reg <= 9'h0;
                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                            if (8'h9e == _T_807) begin
                                                                                                                                                                                                              data_reg <= 9'h0;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                              if (8'h9d == _T_807) begin
                                                                                                                                                                                                                data_reg <= 9'h0;
                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                if (8'h9c == _T_807) begin
                                                                                                                                                                                                                  data_reg <= 9'h0;
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                  if (8'h9b == _T_807) begin
                                                                                                                                                                                                                    data_reg <= 9'h0;
                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                    if (8'h9a == _T_807) begin
                                                                                                                                                                                                                      data_reg <= 9'h0;
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                      if (8'h99 == _T_807) begin
                                                                                                                                                                                                                        data_reg <= 9'h0;
                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                        if (8'h98 == _T_807) begin
                                                                                                                                                                                                                          data_reg <= 9'h0;
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                          if (8'h97 == _T_807) begin
                                                                                                                                                                                                                            data_reg <= 9'h0;
                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                            if (8'h96 == _T_807) begin
                                                                                                                                                                                                                              data_reg <= 9'h0;
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                              if (8'h95 == _T_807) begin
                                                                                                                                                                                                                                data_reg <= 9'h0;
                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                if (8'h94 == _T_807) begin
                                                                                                                                                                                                                                  data_reg <= 9'h0;
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                  if (8'h93 == _T_807) begin
                                                                                                                                                                                                                                    data_reg <= 9'h0;
                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                    if (8'h92 == _T_807) begin
                                                                                                                                                                                                                                      data_reg <= 9'h0;
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                      if (8'h91 == _T_807) begin
                                                                                                                                                                                                                                        data_reg <= 9'h0;
                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                        if (8'h90 == _T_807) begin
                                                                                                                                                                                                                                          data_reg <= 9'h0;
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                          if (8'h8f == _T_807) begin
                                                                                                                                                                                                                                            data_reg <= 9'h0;
                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                            if (8'h8e == _T_807) begin
                                                                                                                                                                                                                                              data_reg <= 9'h0;
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                              if (8'h8d == _T_807) begin
                                                                                                                                                                                                                                                data_reg <= 9'h0;
                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                if (8'h8c == _T_807) begin
                                                                                                                                                                                                                                                  data_reg <= 9'h0;
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                  if (8'h8b == _T_807) begin
                                                                                                                                                                                                                                                    data_reg <= 9'h0;
                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                    if (8'h8a == _T_807) begin
                                                                                                                                                                                                                                                      data_reg <= 9'h0;
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                      if (8'h89 == _T_807) begin
                                                                                                                                                                                                                                                        data_reg <= 9'h0;
                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                        if (8'h88 == _T_807) begin
                                                                                                                                                                                                                                                          data_reg <= 9'h0;
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                          if (8'h87 == _T_807) begin
                                                                                                                                                                                                                                                            data_reg <= 9'h0;
                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                            if (8'h86 == _T_807) begin
                                                                                                                                                                                                                                                              data_reg <= 9'h0;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                              if (8'h85 == _T_807) begin
                                                                                                                                                                                                                                                                data_reg <= 9'h0;
                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                if (8'h84 == _T_807) begin
                                                                                                                                                                                                                                                                  data_reg <= 9'h0;
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                  if (8'h83 == _T_807) begin
                                                                                                                                                                                                                                                                    data_reg <= 9'h0;
                                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                                    if (8'h82 == _T_807) begin
                                                                                                                                                                                                                                                                      data_reg <= 9'h0;
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                      if (8'h81 == _T_807) begin
                                                                                                                                                                                                                                                                        data_reg <= 9'h0;
                                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                                        if (8'h80 == _T_807) begin
                                                                                                                                                                                                                                                                          data_reg <= 9'h0;
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                          if (8'h7f == _T_807) begin
                                                                                                                                                                                                                                                                            data_reg <= 9'h0;
                                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                                            if (8'h7e == _T_807) begin
                                                                                                                                                                                                                                                                              data_reg <= 9'h0;
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                              if (8'h7d == _T_807) begin
                                                                                                                                                                                                                                                                                data_reg <= 9'h0;
                                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                                if (8'h7c == _T_807) begin
                                                                                                                                                                                                                                                                                  data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                  if (8'h7b == _T_807) begin
                                                                                                                                                                                                                                                                                    data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                                                    if (8'h7a == _T_807) begin
                                                                                                                                                                                                                                                                                      data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                      if (8'h79 == _T_807) begin
                                                                                                                                                                                                                                                                                        data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                                                        if (8'h78 == _T_807) begin
                                                                                                                                                                                                                                                                                          data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                          if (8'h77 == _T_807) begin
                                                                                                                                                                                                                                                                                            data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                                                            if (8'h76 == _T_807) begin
                                                                                                                                                                                                                                                                                              data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                              if (8'h75 == _T_807) begin
                                                                                                                                                                                                                                                                                                data_reg <= 9'h116;
                                                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                                                if (8'h74 == _T_807) begin
                                                                                                                                                                                                                                                                                                  data_reg <= 9'h102;
                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                  if (8'h73 == _T_807) begin
                                                                                                                                                                                                                                                                                                    data_reg <= 9'h101;
                                                                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                                                                    if (8'h72 == _T_807) begin
                                                                                                                                                                                                                                                                                                      data_reg <= 9'h78;
                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                      if (8'h71 == _T_807) begin
                                                                                                                                                                                                                                                                                                        data_reg <= 9'h73;
                                                                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                                                                        if (8'h70 == _T_807) begin
                                                                                                                                                                                                                                                                                                          data_reg <= 9'h72;
                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                          if (8'h6f == _T_807) begin
                                                                                                                                                                                                                                                                                                            data_reg <= 9'h6f;
                                                                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                                                                            if (8'h6e == _T_807) begin
                                                                                                                                                                                                                                                                                                              data_reg <= 9'h6d;
                                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                              if (8'h6d == _T_807) begin
                                                                                                                                                                                                                                                                                                                data_reg <= 9'h66;
                                                                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                                                                if (8'h6c == _T_807) begin
                                                                                                                                                                                                                                                                                                                  data_reg <= 9'h61;
                                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                                  if (8'h6b == _T_807) begin
                                                                                                                                                                                                                                                                                                                    data_reg <= 9'h35;
                                                                                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                                                                                    if (8'h6a == _T_807) begin
                                                                                                                                                                                                                                                                                                                      data_reg <= 9'h32;
                                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                                      if (8'h69 == _T_807) begin
                                                                                                                                                                                                                                                                                                                        data_reg <= 9'h30;
                                                                                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                                                                                        if (8'h68 == _T_807) begin
                                                                                                                                                                                                                                                                                                                          data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                                          if (8'h67 == _T_807) begin
                                                                                                                                                                                                                                                                                                                            data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                                                                                            if (8'h66 == _T_807) begin
                                                                                                                                                                                                                                                                                                                              data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                                              if (8'h65 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                                                                                if (8'h64 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                  data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                                                  if (8'h63 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                    data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                                                                                                    if (8'h62 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                      data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                                                      if (8'h61 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                        data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                                                                                                        if (8'h60 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                          data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                                                          if (8'h5f == _T_807) begin
                                                                                                                                                                                                                                                                                                                                            data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                                                                                                            if (8'h5e == _T_807) begin
                                                                                                                                                                                                                                                                                                                                              data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                                                              if (8'h5d == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                                                                                                if (8'h5c == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                  data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                                                                  if (8'h5b == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                    data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                                                                                                                    if (8'h5a == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                      data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                                                                      if (8'h59 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                        data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                                                                                                                        if (8'h58 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                          data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                                                                          if (8'h57 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                            data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                                                                                                                            if (8'h56 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                              data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                                                                              if (8'h55 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                                                                                                                if (8'h54 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                  data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                                                                                  if (8'h53 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                    data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                                                                                                                                    if (8'h52 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                      data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                                                                                      if (8'h51 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                        data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                                                                                                                                        if (8'h50 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                          data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                                                                                          if (8'h4f == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                            data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                                                                                                                                            if (8'h4e == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                              data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                                                                                              if (8'h4d == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                                                                                                                                if (8'h4c == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                  data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                                                                                                  if (8'h4b == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                    data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                                                                                                                                                    if (8'h4a == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                      data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                                                                                                      if (8'h49 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                        data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                                                                                                                                                        if (8'h48 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                          data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                                                                                                          if (8'h47 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                            data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                                                                                                                                                            if (8'h46 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                              data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                                                                                                              if (8'h45 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                                                                                                                                                if (8'h44 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                  data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                                                                                                                  if (8'h43 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                    data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                                                                                                                                                                    if (8'h42 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                      data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                                                                                                                      if (8'h41 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                        data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                                                                                                                                                                        if (8'h40 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                          data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                                                                                                                          if (8'h3f == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                            data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                                                                                                                                                                            if (8'h3e == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                              data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                                                                                                                              if (8'h3d == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                if (8'h3c == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                  data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                  if (8'h3b == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                    data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                    if (8'h3a == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                      data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                      if (8'h39 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                        data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                        if (8'h38 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                          data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                          if (8'h37 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                            data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                            if (8'h36 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                              data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                              if (8'h35 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                if (8'h34 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                  data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                  if (8'h33 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                    data_reg <= 9'h6c;
                                                                                                                                                                                                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                    if (8'h32 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                      data_reg <= 9'h69;
                                                                                                                                                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                      if (8'h31 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                        data_reg <= 9'h65;
                                                                                                                                                                                                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                        if (8'h30 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                          data_reg <= 9'h36;
                                                                                                                                                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                          if (8'h2f == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                            data_reg <= 9'h34;
                                                                                                                                                                                                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                            if (8'h2e == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                              data_reg <= 9'h33;
                                                                                                                                                                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                              if (8'h2d == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                data_reg <= 9'h31;
                                                                                                                                                                                                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                if (8'h2c == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                  data_reg <= 9'ha;
                                                                                                                                                                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                  if (8'h2b == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                    data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                    if (8'h2a == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                      data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                      if (8'h29 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                        data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                        if (8'h28 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                          data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                          if (8'h27 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                            data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                            if (8'h26 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                              data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                              if (8'h25 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                if (8'h24 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                  data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                  if (8'h23 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    if (8'h22 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                      data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                      if (8'h21 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                        data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                        if (8'h20 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                          data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                          if (8'h1f == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                            data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                            if (8'h1e == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              if (8'h1d == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                if (8'h1c == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  if (8'h1b == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    if (8'h1a == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      if (8'h19 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        if (8'h18 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          if (8'h17 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            if (8'h16 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              if (8'h15 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                if (8'h14 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  data_reg <= 9'h74;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  if (8'h13 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    data_reg <= 9'h20;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    if (8'h12 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      if (8'h11 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        if (8'h10 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          if (8'hf == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            if (8'he == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              if (8'hd == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                if (8'hc == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  if (8'hb == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    if (8'ha == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      if (8'h9 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        if (8'h8 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          if (8'h7 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            if (8'h6 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              if (8'h5 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                if (8'h4 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  if (8'h3 == _T_807) begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    data_reg <= 9'h11d;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    data_reg <= 9'h0;
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                              end
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                          end
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                      end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                  end
                                                                                                                                                                                                                end
                                                                                                                                                                                                              end
                                                                                                                                                                                                            end
                                                                                                                                                                                                          end
                                                                                                                                                                                                        end
                                                                                                                                                                                                      end
                                                                                                                                                                                                    end
                                                                                                                                                                                                  end
                                                                                                                                                                                                end
                                                                                                                                                                                              end
                                                                                                                                                                                            end
                                                                                                                                                                                          end
                                                                                                                                                                                        end
                                                                                                                                                                                      end
                                                                                                                                                                                    end
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end
                                                                                                                                                                  end
                                                                                                                                                                end
                                                                                                                                                              end
                                                                                                                                                            end
                                                                                                                                                          end
                                                                                                                                                        end
                                                                                                                                                      end
                                                                                                                                                    end
                                                                                                                                                  end
                                                                                                                                                end
                                                                                                                                              end
                                                                                                                                            end
                                                                                                                                          end
                                                                                                                                        end
                                                                                                                                      end
                                                                                                                                    end
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_1551 & _T_797) begin
          $fwrite(32'h80000002,"DEC ERR\n"); // @[GunzipHuffDecoder.scala 54:13:@551.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module GunzipLenDistLut( // @[:@579.2]
  input         clock, // @[:@580.4]
  input         reset, // @[:@581.4]
  input         io_data_in_valid, // @[:@582.4]
  output        io_data_in_ready, // @[:@582.4]
  input         io_data_in_bits, // @[:@582.4]
  input         io_enable, // @[:@582.4]
  input  [8:0]  io_lut_idx, // @[:@582.4]
  output        io_done, // @[:@582.4]
  output [14:0] io_lut_out // @[:@582.4]
);
  reg [1:0] state; // @[GunzipLenDistLut.scala 66:22:@644.4]
  reg [31:0] _RAND_0;
  reg  done_reg; // @[GunzipLenDistLut.scala 69:21:@645.4]
  reg [31:0] _RAND_1;
  reg [14:0] out_reg; // @[GunzipLenDistLut.scala 70:20:@646.4]
  reg [31:0] _RAND_2;
  reg [8:0] val_init; // @[GunzipLenDistLut.scala 75:22:@649.4]
  reg [31:0] _RAND_3;
  reg [4:0] ext_idx; // @[GunzipLenDistLut.scala 76:21:@650.4]
  reg [31:0] _RAND_4;
  reg [4:0] ext_lim; // @[GunzipLenDistLut.scala 77:21:@651.4]
  reg [31:0] _RAND_5;
  reg [6:0] ext_val; // @[GunzipLenDistLut.scala 78:21:@652.4]
  reg [31:0] _RAND_6;
  wire  _T_154; // @[Conditional.scala 37:30:@653.4]
  wire  _T_156; // @[GunzipLenDistLut.scala 82:26:@655.6]
  wire  _T_157; // @[GunzipLenDistLut.scala 82:23:@656.6]
  wire [4:0] _T_159; // @[:@658.8]
  wire [14:0] _GEN_8; // @[GunzipLenDistLut.scala 83:32:@659.8]
  wire [14:0] _GEN_9; // @[GunzipLenDistLut.scala 83:32:@659.8]
  wire [14:0] _GEN_10; // @[GunzipLenDistLut.scala 83:32:@659.8]
  wire [14:0] _GEN_11; // @[GunzipLenDistLut.scala 83:32:@659.8]
  wire [14:0] _GEN_12; // @[GunzipLenDistLut.scala 83:32:@659.8]
  wire [14:0] _GEN_13; // @[GunzipLenDistLut.scala 83:32:@659.8]
  wire [14:0] _GEN_14; // @[GunzipLenDistLut.scala 83:32:@659.8]
  wire [14:0] _GEN_15; // @[GunzipLenDistLut.scala 83:32:@659.8]
  wire [14:0] _GEN_16; // @[GunzipLenDistLut.scala 83:32:@659.8]
  wire [14:0] _GEN_17; // @[GunzipLenDistLut.scala 83:32:@659.8]
  wire [14:0] _GEN_18; // @[GunzipLenDistLut.scala 83:32:@659.8]
  wire [14:0] _GEN_19; // @[GunzipLenDistLut.scala 83:32:@659.8]
  wire [14:0] _GEN_20; // @[GunzipLenDistLut.scala 83:32:@659.8]
  wire [14:0] _GEN_21; // @[GunzipLenDistLut.scala 83:32:@659.8]
  wire [14:0] _GEN_22; // @[GunzipLenDistLut.scala 83:32:@659.8]
  wire [14:0] _GEN_23; // @[GunzipLenDistLut.scala 83:32:@659.8]
  wire [14:0] _GEN_24; // @[GunzipLenDistLut.scala 83:32:@659.8]
  wire [14:0] _GEN_25; // @[GunzipLenDistLut.scala 83:32:@659.8]
  wire [14:0] _GEN_26; // @[GunzipLenDistLut.scala 83:32:@659.8]
  wire [14:0] _GEN_27; // @[GunzipLenDistLut.scala 83:32:@659.8]
  wire [14:0] _GEN_28; // @[GunzipLenDistLut.scala 83:32:@659.8]
  wire  _T_161; // @[GunzipLenDistLut.scala 83:32:@659.8]
  wire [14:0] _GEN_30; // @[GunzipLenDistLut.scala 85:20:@663.10]
  wire [14:0] _GEN_31; // @[GunzipLenDistLut.scala 85:20:@663.10]
  wire [14:0] _GEN_32; // @[GunzipLenDistLut.scala 85:20:@663.10]
  wire [14:0] _GEN_33; // @[GunzipLenDistLut.scala 85:20:@663.10]
  wire [14:0] _GEN_34; // @[GunzipLenDistLut.scala 85:20:@663.10]
  wire [14:0] _GEN_35; // @[GunzipLenDistLut.scala 85:20:@663.10]
  wire [14:0] _GEN_36; // @[GunzipLenDistLut.scala 85:20:@663.10]
  wire [14:0] _GEN_37; // @[GunzipLenDistLut.scala 85:20:@663.10]
  wire [14:0] _GEN_38; // @[GunzipLenDistLut.scala 85:20:@663.10]
  wire [14:0] _GEN_39; // @[GunzipLenDistLut.scala 85:20:@663.10]
  wire [14:0] _GEN_40; // @[GunzipLenDistLut.scala 85:20:@663.10]
  wire [14:0] _GEN_41; // @[GunzipLenDistLut.scala 85:20:@663.10]
  wire [14:0] _GEN_42; // @[GunzipLenDistLut.scala 85:20:@663.10]
  wire [14:0] _GEN_43; // @[GunzipLenDistLut.scala 85:20:@663.10]
  wire [14:0] _GEN_44; // @[GunzipLenDistLut.scala 85:20:@663.10]
  wire [14:0] _GEN_45; // @[GunzipLenDistLut.scala 85:20:@663.10]
  wire [14:0] _GEN_46; // @[GunzipLenDistLut.scala 85:20:@663.10]
  wire [14:0] _GEN_47; // @[GunzipLenDistLut.scala 85:20:@663.10]
  wire [14:0] _GEN_48; // @[GunzipLenDistLut.scala 85:20:@663.10]
  wire [14:0] _GEN_49; // @[GunzipLenDistLut.scala 85:20:@663.10]
  wire [14:0] _GEN_50; // @[GunzipLenDistLut.scala 85:20:@663.10]
  wire [14:0] _GEN_51; // @[GunzipLenDistLut.scala 85:20:@663.10]
  wire [14:0] _GEN_52; // @[GunzipLenDistLut.scala 85:20:@663.10]
  wire [14:0] _GEN_53; // @[GunzipLenDistLut.scala 85:20:@663.10]
  wire [14:0] _GEN_54; // @[GunzipLenDistLut.scala 85:20:@663.10]
  wire [14:0] _GEN_55; // @[GunzipLenDistLut.scala 85:20:@663.10]
  wire [14:0] _GEN_56; // @[GunzipLenDistLut.scala 85:20:@663.10]
  wire [14:0] _GEN_57; // @[GunzipLenDistLut.scala 85:20:@663.10]
  wire [15:0] _T_168; // @[GunzipLenDistLut.scala 87:39:@666.10]
  wire [15:0] _T_169; // @[GunzipLenDistLut.scala 87:39:@667.10]
  wire [14:0] _T_170; // @[GunzipLenDistLut.scala 87:39:@668.10]
  wire [1:0] _GEN_116; // @[GunzipLenDistLut.scala 83:39:@660.8]
  wire [14:0] _GEN_117; // @[GunzipLenDistLut.scala 83:39:@660.8]
  wire [4:0] _GEN_118; // @[GunzipLenDistLut.scala 83:39:@660.8]
  wire [14:0] _GEN_119; // @[GunzipLenDistLut.scala 83:39:@660.8]
  wire [6:0] _GEN_120; // @[GunzipLenDistLut.scala 83:39:@660.8]
  wire  _GEN_121; // @[GunzipLenDistLut.scala 83:39:@660.8]
  wire [14:0] _GEN_122; // @[GunzipLenDistLut.scala 83:39:@660.8]
  wire [1:0] _GEN_123; // @[GunzipLenDistLut.scala 82:36:@657.6]
  wire [14:0] _GEN_124; // @[GunzipLenDistLut.scala 82:36:@657.6]
  wire [4:0] _GEN_125; // @[GunzipLenDistLut.scala 82:36:@657.6]
  wire [14:0] _GEN_126; // @[GunzipLenDistLut.scala 82:36:@657.6]
  wire [6:0] _GEN_127; // @[GunzipLenDistLut.scala 82:36:@657.6]
  wire  _GEN_128; // @[GunzipLenDistLut.scala 82:36:@657.6]
  wire [14:0] _GEN_129; // @[GunzipLenDistLut.scala 82:36:@657.6]
  wire  _T_175; // @[Conditional.scala 37:30:@681.6]
  wire  _T_181; // @[Conditional.scala 37:30:@687.10]
  wire [5:0] _T_182; // @[GunzipLenDistLut.scala 50:33:@689.12]
  wire [6:0] _T_183; // @[Cat.scala 30:58:@690.12]
  wire  _T_185; // @[Conditional.scala 37:30:@694.12]
  wire [4:0] _T_186; // @[GunzipLenDistLut.scala 51:33:@696.14]
  wire  _T_187; // @[GunzipLenDistLut.scala 51:70:@697.14]
  wire [6:0] _T_189; // @[Cat.scala 30:58:@699.14]
  wire  _T_191; // @[Conditional.scala 37:30:@703.14]
  wire [3:0] _T_192; // @[GunzipLenDistLut.scala 52:33:@705.16]
  wire [1:0] _T_193; // @[GunzipLenDistLut.scala 52:70:@706.16]
  wire [6:0] _T_195; // @[Cat.scala 30:58:@708.16]
  wire  _T_197; // @[Conditional.scala 37:30:@712.16]
  wire [2:0] _T_198; // @[GunzipLenDistLut.scala 53:33:@714.18]
  wire [2:0] _T_199; // @[GunzipLenDistLut.scala 53:70:@715.18]
  wire [6:0] _T_201; // @[Cat.scala 30:58:@717.18]
  wire  _T_203; // @[Conditional.scala 37:30:@721.18]
  wire [1:0] _T_204; // @[GunzipLenDistLut.scala 54:33:@723.20]
  wire [3:0] _T_205; // @[GunzipLenDistLut.scala 54:70:@724.20]
  wire [6:0] _T_207; // @[Cat.scala 30:58:@726.20]
  wire  _T_209; // @[Conditional.scala 37:30:@730.20]
  wire  _T_210; // @[GunzipLenDistLut.scala 55:33:@732.22]
  wire [4:0] _T_211; // @[GunzipLenDistLut.scala 55:70:@733.22]
  wire [6:0] _T_213; // @[Cat.scala 30:58:@735.22]
  wire [6:0] _GEN_130; // @[Conditional.scala 39:67:@731.20]
  wire [6:0] _GEN_131; // @[Conditional.scala 39:67:@722.18]
  wire [6:0] _GEN_132; // @[Conditional.scala 39:67:@713.16]
  wire [6:0] _GEN_133; // @[Conditional.scala 39:67:@704.14]
  wire [6:0] _GEN_134; // @[Conditional.scala 39:67:@695.12]
  wire [6:0] _GEN_135; // @[Conditional.scala 40:58:@688.10]
  wire [5:0] _T_215; // @[GunzipLenDistLut.scala 100:28:@739.10]
  wire [4:0] _T_216; // @[GunzipLenDistLut.scala 100:28:@740.10]
  wire  _T_217; // @[GunzipLenDistLut.scala 102:22:@742.10]
  wire [1:0] _GEN_136; // @[GunzipLenDistLut.scala 102:35:@743.10]
  wire [6:0] _GEN_138; // @[GunzipLenDistLut.scala 97:31:@683.8]
  wire [4:0] _GEN_139; // @[GunzipLenDistLut.scala 97:31:@683.8]
  wire [1:0] _GEN_140; // @[GunzipLenDistLut.scala 97:31:@683.8]
  wire  _T_218; // @[Conditional.scala 37:30:@749.8]
  wire [8:0] _GEN_159; // @[GunzipLenDistLut.scala 110:27:@753.10]
  wire [9:0] _T_220; // @[GunzipLenDistLut.scala 110:27:@753.10]
  wire [8:0] _T_221; // @[GunzipLenDistLut.scala 110:27:@754.10]
  wire [1:0] _GEN_141; // @[Conditional.scala 39:67:@750.8]
  wire [14:0] _GEN_143; // @[Conditional.scala 39:67:@750.8]
  wire  _GEN_144; // @[Conditional.scala 39:67:@682.6]
  wire [6:0] _GEN_145; // @[Conditional.scala 39:67:@682.6]
  wire [4:0] _GEN_146; // @[Conditional.scala 39:67:@682.6]
  wire [1:0] _GEN_147; // @[Conditional.scala 39:67:@682.6]
  wire  _GEN_148; // @[Conditional.scala 39:67:@682.6]
  wire [14:0] _GEN_149; // @[Conditional.scala 39:67:@682.6]
  wire [1:0] _GEN_150; // @[Conditional.scala 40:58:@654.4]
  wire [14:0] _GEN_151; // @[Conditional.scala 40:58:@654.4]
  wire [14:0] _GEN_153; // @[Conditional.scala 40:58:@654.4]
  wire  _GEN_157; // @[Conditional.scala 40:58:@654.4]
  assign _T_154 = 2'h0 == state; // @[Conditional.scala 37:30:@653.4]
  assign _T_156 = io_done == 1'h0; // @[GunzipLenDistLut.scala 82:26:@655.6]
  assign _T_157 = io_enable & _T_156; // @[GunzipLenDistLut.scala 82:23:@656.6]
  assign _T_159 = io_lut_idx[4:0]; // @[:@658.8]
  assign _GEN_8 = 5'h8 == _T_159 ? 15'h1 : 15'h0; // @[GunzipLenDistLut.scala 83:32:@659.8]
  assign _GEN_9 = 5'h9 == _T_159 ? 15'h1 : _GEN_8; // @[GunzipLenDistLut.scala 83:32:@659.8]
  assign _GEN_10 = 5'ha == _T_159 ? 15'h1 : _GEN_9; // @[GunzipLenDistLut.scala 83:32:@659.8]
  assign _GEN_11 = 5'hb == _T_159 ? 15'h1 : _GEN_10; // @[GunzipLenDistLut.scala 83:32:@659.8]
  assign _GEN_12 = 5'hc == _T_159 ? 15'h2 : _GEN_11; // @[GunzipLenDistLut.scala 83:32:@659.8]
  assign _GEN_13 = 5'hd == _T_159 ? 15'h2 : _GEN_12; // @[GunzipLenDistLut.scala 83:32:@659.8]
  assign _GEN_14 = 5'he == _T_159 ? 15'h2 : _GEN_13; // @[GunzipLenDistLut.scala 83:32:@659.8]
  assign _GEN_15 = 5'hf == _T_159 ? 15'h2 : _GEN_14; // @[GunzipLenDistLut.scala 83:32:@659.8]
  assign _GEN_16 = 5'h10 == _T_159 ? 15'h3 : _GEN_15; // @[GunzipLenDistLut.scala 83:32:@659.8]
  assign _GEN_17 = 5'h11 == _T_159 ? 15'h3 : _GEN_16; // @[GunzipLenDistLut.scala 83:32:@659.8]
  assign _GEN_18 = 5'h12 == _T_159 ? 15'h3 : _GEN_17; // @[GunzipLenDistLut.scala 83:32:@659.8]
  assign _GEN_19 = 5'h13 == _T_159 ? 15'h3 : _GEN_18; // @[GunzipLenDistLut.scala 83:32:@659.8]
  assign _GEN_20 = 5'h14 == _T_159 ? 15'h4 : _GEN_19; // @[GunzipLenDistLut.scala 83:32:@659.8]
  assign _GEN_21 = 5'h15 == _T_159 ? 15'h4 : _GEN_20; // @[GunzipLenDistLut.scala 83:32:@659.8]
  assign _GEN_22 = 5'h16 == _T_159 ? 15'h4 : _GEN_21; // @[GunzipLenDistLut.scala 83:32:@659.8]
  assign _GEN_23 = 5'h17 == _T_159 ? 15'h4 : _GEN_22; // @[GunzipLenDistLut.scala 83:32:@659.8]
  assign _GEN_24 = 5'h18 == _T_159 ? 15'h5 : _GEN_23; // @[GunzipLenDistLut.scala 83:32:@659.8]
  assign _GEN_25 = 5'h19 == _T_159 ? 15'h5 : _GEN_24; // @[GunzipLenDistLut.scala 83:32:@659.8]
  assign _GEN_26 = 5'h1a == _T_159 ? 15'h5 : _GEN_25; // @[GunzipLenDistLut.scala 83:32:@659.8]
  assign _GEN_27 = 5'h1b == _T_159 ? 15'h5 : _GEN_26; // @[GunzipLenDistLut.scala 83:32:@659.8]
  assign _GEN_28 = 5'h1c == _T_159 ? 15'h0 : _GEN_27; // @[GunzipLenDistLut.scala 83:32:@659.8]
  assign _T_161 = _GEN_28 > 15'h0; // @[GunzipLenDistLut.scala 83:32:@659.8]
  assign _GEN_30 = 5'h1 == _T_159 ? 15'h4 : 15'h3; // @[GunzipLenDistLut.scala 85:20:@663.10]
  assign _GEN_31 = 5'h2 == _T_159 ? 15'h5 : _GEN_30; // @[GunzipLenDistLut.scala 85:20:@663.10]
  assign _GEN_32 = 5'h3 == _T_159 ? 15'h6 : _GEN_31; // @[GunzipLenDistLut.scala 85:20:@663.10]
  assign _GEN_33 = 5'h4 == _T_159 ? 15'h7 : _GEN_32; // @[GunzipLenDistLut.scala 85:20:@663.10]
  assign _GEN_34 = 5'h5 == _T_159 ? 15'h8 : _GEN_33; // @[GunzipLenDistLut.scala 85:20:@663.10]
  assign _GEN_35 = 5'h6 == _T_159 ? 15'h9 : _GEN_34; // @[GunzipLenDistLut.scala 85:20:@663.10]
  assign _GEN_36 = 5'h7 == _T_159 ? 15'ha : _GEN_35; // @[GunzipLenDistLut.scala 85:20:@663.10]
  assign _GEN_37 = 5'h8 == _T_159 ? 15'hb : _GEN_36; // @[GunzipLenDistLut.scala 85:20:@663.10]
  assign _GEN_38 = 5'h9 == _T_159 ? 15'hd : _GEN_37; // @[GunzipLenDistLut.scala 85:20:@663.10]
  assign _GEN_39 = 5'ha == _T_159 ? 15'hf : _GEN_38; // @[GunzipLenDistLut.scala 85:20:@663.10]
  assign _GEN_40 = 5'hb == _T_159 ? 15'h11 : _GEN_39; // @[GunzipLenDistLut.scala 85:20:@663.10]
  assign _GEN_41 = 5'hc == _T_159 ? 15'h13 : _GEN_40; // @[GunzipLenDistLut.scala 85:20:@663.10]
  assign _GEN_42 = 5'hd == _T_159 ? 15'h17 : _GEN_41; // @[GunzipLenDistLut.scala 85:20:@663.10]
  assign _GEN_43 = 5'he == _T_159 ? 15'h1b : _GEN_42; // @[GunzipLenDistLut.scala 85:20:@663.10]
  assign _GEN_44 = 5'hf == _T_159 ? 15'h1f : _GEN_43; // @[GunzipLenDistLut.scala 85:20:@663.10]
  assign _GEN_45 = 5'h10 == _T_159 ? 15'h23 : _GEN_44; // @[GunzipLenDistLut.scala 85:20:@663.10]
  assign _GEN_46 = 5'h11 == _T_159 ? 15'h2b : _GEN_45; // @[GunzipLenDistLut.scala 85:20:@663.10]
  assign _GEN_47 = 5'h12 == _T_159 ? 15'h33 : _GEN_46; // @[GunzipLenDistLut.scala 85:20:@663.10]
  assign _GEN_48 = 5'h13 == _T_159 ? 15'h3b : _GEN_47; // @[GunzipLenDistLut.scala 85:20:@663.10]
  assign _GEN_49 = 5'h14 == _T_159 ? 15'h43 : _GEN_48; // @[GunzipLenDistLut.scala 85:20:@663.10]
  assign _GEN_50 = 5'h15 == _T_159 ? 15'h53 : _GEN_49; // @[GunzipLenDistLut.scala 85:20:@663.10]
  assign _GEN_51 = 5'h16 == _T_159 ? 15'h63 : _GEN_50; // @[GunzipLenDistLut.scala 85:20:@663.10]
  assign _GEN_52 = 5'h17 == _T_159 ? 15'h73 : _GEN_51; // @[GunzipLenDistLut.scala 85:20:@663.10]
  assign _GEN_53 = 5'h18 == _T_159 ? 15'h83 : _GEN_52; // @[GunzipLenDistLut.scala 85:20:@663.10]
  assign _GEN_54 = 5'h19 == _T_159 ? 15'ha3 : _GEN_53; // @[GunzipLenDistLut.scala 85:20:@663.10]
  assign _GEN_55 = 5'h1a == _T_159 ? 15'hc3 : _GEN_54; // @[GunzipLenDistLut.scala 85:20:@663.10]
  assign _GEN_56 = 5'h1b == _T_159 ? 15'he3 : _GEN_55; // @[GunzipLenDistLut.scala 85:20:@663.10]
  assign _GEN_57 = 5'h1c == _T_159 ? 15'h102 : _GEN_56; // @[GunzipLenDistLut.scala 85:20:@663.10]
  assign _T_168 = _GEN_28 - 15'h1; // @[GunzipLenDistLut.scala 87:39:@666.10]
  assign _T_169 = $unsigned(_T_168); // @[GunzipLenDistLut.scala 87:39:@667.10]
  assign _T_170 = _T_169[14:0]; // @[GunzipLenDistLut.scala 87:39:@668.10]
  assign _GEN_116 = _T_161 ? 2'h1 : 2'h0; // @[GunzipLenDistLut.scala 83:39:@660.8]
  assign _GEN_117 = _T_161 ? _GEN_57 : {{6'd0}, val_init}; // @[GunzipLenDistLut.scala 83:39:@660.8]
  assign _GEN_118 = _T_161 ? 5'h0 : ext_idx; // @[GunzipLenDistLut.scala 83:39:@660.8]
  assign _GEN_119 = _T_161 ? _T_170 : {{10'd0}, ext_lim}; // @[GunzipLenDistLut.scala 83:39:@660.8]
  assign _GEN_120 = _T_161 ? 7'h0 : ext_val; // @[GunzipLenDistLut.scala 83:39:@660.8]
  assign _GEN_121 = _T_161 ? 1'h0 : 1'h1; // @[GunzipLenDistLut.scala 83:39:@660.8]
  assign _GEN_122 = _T_161 ? out_reg : _GEN_57; // @[GunzipLenDistLut.scala 83:39:@660.8]
  assign _GEN_123 = _T_157 ? _GEN_116 : state; // @[GunzipLenDistLut.scala 82:36:@657.6]
  assign _GEN_124 = _T_157 ? _GEN_117 : {{6'd0}, val_init}; // @[GunzipLenDistLut.scala 82:36:@657.6]
  assign _GEN_125 = _T_157 ? _GEN_118 : ext_idx; // @[GunzipLenDistLut.scala 82:36:@657.6]
  assign _GEN_126 = _T_157 ? _GEN_119 : {{10'd0}, ext_lim}; // @[GunzipLenDistLut.scala 82:36:@657.6]
  assign _GEN_127 = _T_157 ? _GEN_120 : ext_val; // @[GunzipLenDistLut.scala 82:36:@657.6]
  assign _GEN_128 = _T_157 ? _GEN_121 : 1'h0; // @[GunzipLenDistLut.scala 82:36:@657.6]
  assign _GEN_129 = _T_157 ? _GEN_122 : out_reg; // @[GunzipLenDistLut.scala 82:36:@657.6]
  assign _T_175 = 2'h1 == state; // @[Conditional.scala 37:30:@681.6]
  assign _T_181 = 5'h0 == ext_idx; // @[Conditional.scala 37:30:@687.10]
  assign _T_182 = ext_val[6:1]; // @[GunzipLenDistLut.scala 50:33:@689.12]
  assign _T_183 = {_T_182,io_data_in_bits}; // @[Cat.scala 30:58:@690.12]
  assign _T_185 = 5'h1 == ext_idx; // @[Conditional.scala 37:30:@694.12]
  assign _T_186 = ext_val[6:2]; // @[GunzipLenDistLut.scala 51:33:@696.14]
  assign _T_187 = ext_val[0]; // @[GunzipLenDistLut.scala 51:70:@697.14]
  assign _T_189 = {_T_186,io_data_in_bits,_T_187}; // @[Cat.scala 30:58:@699.14]
  assign _T_191 = 5'h2 == ext_idx; // @[Conditional.scala 37:30:@703.14]
  assign _T_192 = ext_val[6:3]; // @[GunzipLenDistLut.scala 52:33:@705.16]
  assign _T_193 = ext_val[1:0]; // @[GunzipLenDistLut.scala 52:70:@706.16]
  assign _T_195 = {_T_192,io_data_in_bits,_T_193}; // @[Cat.scala 30:58:@708.16]
  assign _T_197 = 5'h3 == ext_idx; // @[Conditional.scala 37:30:@712.16]
  assign _T_198 = ext_val[6:4]; // @[GunzipLenDistLut.scala 53:33:@714.18]
  assign _T_199 = ext_val[2:0]; // @[GunzipLenDistLut.scala 53:70:@715.18]
  assign _T_201 = {_T_198,io_data_in_bits,_T_199}; // @[Cat.scala 30:58:@717.18]
  assign _T_203 = 5'h4 == ext_idx; // @[Conditional.scala 37:30:@721.18]
  assign _T_204 = ext_val[6:5]; // @[GunzipLenDistLut.scala 54:33:@723.20]
  assign _T_205 = ext_val[3:0]; // @[GunzipLenDistLut.scala 54:70:@724.20]
  assign _T_207 = {_T_204,io_data_in_bits,_T_205}; // @[Cat.scala 30:58:@726.20]
  assign _T_209 = 5'h5 == ext_idx; // @[Conditional.scala 37:30:@730.20]
  assign _T_210 = ext_val[6]; // @[GunzipLenDistLut.scala 55:33:@732.22]
  assign _T_211 = ext_val[4:0]; // @[GunzipLenDistLut.scala 55:70:@733.22]
  assign _T_213 = {_T_210,io_data_in_bits,_T_211}; // @[Cat.scala 30:58:@735.22]
  assign _GEN_130 = _T_209 ? _T_213 : 7'h0; // @[Conditional.scala 39:67:@731.20]
  assign _GEN_131 = _T_203 ? _T_207 : _GEN_130; // @[Conditional.scala 39:67:@722.18]
  assign _GEN_132 = _T_197 ? _T_201 : _GEN_131; // @[Conditional.scala 39:67:@713.16]
  assign _GEN_133 = _T_191 ? _T_195 : _GEN_132; // @[Conditional.scala 39:67:@704.14]
  assign _GEN_134 = _T_185 ? _T_189 : _GEN_133; // @[Conditional.scala 39:67:@695.12]
  assign _GEN_135 = _T_181 ? _T_183 : _GEN_134; // @[Conditional.scala 40:58:@688.10]
  assign _T_215 = ext_idx + 5'h1; // @[GunzipLenDistLut.scala 100:28:@739.10]
  assign _T_216 = ext_idx + 5'h1; // @[GunzipLenDistLut.scala 100:28:@740.10]
  assign _T_217 = ext_idx == ext_lim; // @[GunzipLenDistLut.scala 102:22:@742.10]
  assign _GEN_136 = _T_217 ? 2'h2 : state; // @[GunzipLenDistLut.scala 102:35:@743.10]
  assign _GEN_138 = io_data_in_valid ? _GEN_135 : ext_val; // @[GunzipLenDistLut.scala 97:31:@683.8]
  assign _GEN_139 = io_data_in_valid ? _T_216 : ext_idx; // @[GunzipLenDistLut.scala 97:31:@683.8]
  assign _GEN_140 = io_data_in_valid ? _GEN_136 : state; // @[GunzipLenDistLut.scala 97:31:@683.8]
  assign _T_218 = 2'h2 == state; // @[Conditional.scala 37:30:@749.8]
  assign _GEN_159 = {{2'd0}, ext_val}; // @[GunzipLenDistLut.scala 110:27:@753.10]
  assign _T_220 = val_init + _GEN_159; // @[GunzipLenDistLut.scala 110:27:@753.10]
  assign _T_221 = val_init + _GEN_159; // @[GunzipLenDistLut.scala 110:27:@754.10]
  assign _GEN_141 = _T_218 ? 2'h0 : state; // @[Conditional.scala 39:67:@750.8]
  assign _GEN_143 = _T_218 ? {{6'd0}, _T_221} : out_reg; // @[Conditional.scala 39:67:@750.8]
  assign _GEN_144 = _T_175 ? io_data_in_valid : 1'h0; // @[Conditional.scala 39:67:@682.6]
  assign _GEN_145 = _T_175 ? _GEN_138 : ext_val; // @[Conditional.scala 39:67:@682.6]
  assign _GEN_146 = _T_175 ? _GEN_139 : ext_idx; // @[Conditional.scala 39:67:@682.6]
  assign _GEN_147 = _T_175 ? _GEN_140 : _GEN_141; // @[Conditional.scala 39:67:@682.6]
  assign _GEN_148 = _T_175 ? 1'h0 : _T_218; // @[Conditional.scala 39:67:@682.6]
  assign _GEN_149 = _T_175 ? out_reg : _GEN_143; // @[Conditional.scala 39:67:@682.6]
  assign _GEN_150 = _T_154 ? _GEN_123 : _GEN_147; // @[Conditional.scala 40:58:@654.4]
  assign _GEN_151 = _T_154 ? _GEN_124 : {{6'd0}, val_init}; // @[Conditional.scala 40:58:@654.4]
  assign _GEN_153 = _T_154 ? _GEN_126 : {{10'd0}, ext_lim}; // @[Conditional.scala 40:58:@654.4]
  assign _GEN_157 = _T_154 ? 1'h0 : _GEN_144; // @[Conditional.scala 40:58:@654.4]
  assign io_data_in_ready = done_reg ? 1'h0 : _GEN_157; // @[GunzipLenDistLut.scala 72:20:@648.4 GunzipLenDistLut.scala 98:26:@684.10 GunzipLenDistLut.scala 118:22:@760.6]
  assign io_done = done_reg; // @[GunzipLenDistLut.scala 115:11:@758.4]
  assign io_lut_out = out_reg; // @[GunzipLenDistLut.scala 114:14:@757.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  done_reg = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_reg = _RAND_2[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  val_init = _RAND_3[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  ext_idx = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  ext_lim = _RAND_5[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  ext_val = _RAND_6[6:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_154) begin
        if (_T_157) begin
          if (_T_161) begin
            state <= 2'h1;
          end else begin
            state <= 2'h0;
          end
        end
      end else begin
        if (_T_175) begin
          if (io_data_in_valid) begin
            if (_T_217) begin
              state <= 2'h2;
            end
          end
        end else begin
          if (_T_218) begin
            state <= 2'h0;
          end
        end
      end
    end
    if (_T_154) begin
      if (_T_157) begin
        if (_T_161) begin
          done_reg <= 1'h0;
        end else begin
          done_reg <= 1'h1;
        end
      end else begin
        done_reg <= 1'h0;
      end
    end else begin
      if (_T_175) begin
        done_reg <= 1'h0;
      end else begin
        done_reg <= _T_218;
      end
    end
    if (_T_154) begin
      if (_T_157) begin
        if (!(_T_161)) begin
          if (5'h1c == _T_159) begin
            out_reg <= 15'h102;
          end else begin
            if (5'h1b == _T_159) begin
              out_reg <= 15'he3;
            end else begin
              if (5'h1a == _T_159) begin
                out_reg <= 15'hc3;
              end else begin
                if (5'h19 == _T_159) begin
                  out_reg <= 15'ha3;
                end else begin
                  if (5'h18 == _T_159) begin
                    out_reg <= 15'h83;
                  end else begin
                    if (5'h17 == _T_159) begin
                      out_reg <= 15'h73;
                    end else begin
                      if (5'h16 == _T_159) begin
                        out_reg <= 15'h63;
                      end else begin
                        if (5'h15 == _T_159) begin
                          out_reg <= 15'h53;
                        end else begin
                          if (5'h14 == _T_159) begin
                            out_reg <= 15'h43;
                          end else begin
                            if (5'h13 == _T_159) begin
                              out_reg <= 15'h3b;
                            end else begin
                              if (5'h12 == _T_159) begin
                                out_reg <= 15'h33;
                              end else begin
                                if (5'h11 == _T_159) begin
                                  out_reg <= 15'h2b;
                                end else begin
                                  if (5'h10 == _T_159) begin
                                    out_reg <= 15'h23;
                                  end else begin
                                    if (5'hf == _T_159) begin
                                      out_reg <= 15'h1f;
                                    end else begin
                                      if (5'he == _T_159) begin
                                        out_reg <= 15'h1b;
                                      end else begin
                                        if (5'hd == _T_159) begin
                                          out_reg <= 15'h17;
                                        end else begin
                                          if (5'hc == _T_159) begin
                                            out_reg <= 15'h13;
                                          end else begin
                                            if (5'hb == _T_159) begin
                                              out_reg <= 15'h11;
                                            end else begin
                                              if (5'ha == _T_159) begin
                                                out_reg <= 15'hf;
                                              end else begin
                                                if (5'h9 == _T_159) begin
                                                  out_reg <= 15'hd;
                                                end else begin
                                                  if (5'h8 == _T_159) begin
                                                    out_reg <= 15'hb;
                                                  end else begin
                                                    if (5'h7 == _T_159) begin
                                                      out_reg <= 15'ha;
                                                    end else begin
                                                      if (5'h6 == _T_159) begin
                                                        out_reg <= 15'h9;
                                                      end else begin
                                                        if (5'h5 == _T_159) begin
                                                          out_reg <= 15'h8;
                                                        end else begin
                                                          if (5'h4 == _T_159) begin
                                                            out_reg <= 15'h7;
                                                          end else begin
                                                            if (5'h3 == _T_159) begin
                                                              out_reg <= 15'h6;
                                                            end else begin
                                                              if (5'h2 == _T_159) begin
                                                                out_reg <= 15'h5;
                                                              end else begin
                                                                if (5'h1 == _T_159) begin
                                                                  out_reg <= 15'h4;
                                                                end else begin
                                                                  out_reg <= 15'h3;
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (!(_T_175)) begin
        if (_T_218) begin
          out_reg <= {{6'd0}, _T_221};
        end
      end
    end
    val_init <= _GEN_151[8:0];
    if (_T_154) begin
      if (_T_157) begin
        if (_T_161) begin
          ext_idx <= 5'h0;
        end
      end
    end else begin
      if (_T_175) begin
        if (io_data_in_valid) begin
          ext_idx <= _T_216;
        end
      end
    end
    ext_lim <= _GEN_153[4:0];
    if (_T_154) begin
      if (_T_157) begin
        if (_T_161) begin
          ext_val <= 7'h0;
        end
      end
    end else begin
      if (_T_175) begin
        if (io_data_in_valid) begin
          if (_T_181) begin
            ext_val <= _T_183;
          end else begin
            if (_T_185) begin
              ext_val <= _T_189;
            end else begin
              if (_T_191) begin
                ext_val <= _T_195;
              end else begin
                if (_T_197) begin
                  ext_val <= _T_201;
                end else begin
                  if (_T_203) begin
                    ext_val <= _T_207;
                  end else begin
                    if (_T_209) begin
                      ext_val <= _T_213;
                    end else begin
                      ext_val <= 7'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
  end
endmodule
module GunzipHuffDecoder_1( // @[:@763.2]
  input        clock, // @[:@764.4]
  input        reset, // @[:@765.4]
  input        io_data_in_valid, // @[:@766.4]
  output       io_data_in_ready, // @[:@766.4]
  input        io_data_in_bits, // @[:@766.4]
  input        io_enable, // @[:@766.4]
  output [8:0] io_data, // @[:@766.4]
  output       io_valid // @[:@766.4]
);
  reg [8:0] lit_idx; // @[GunzipHuffDecoder.scala 41:24:@768.4]
  reg [31:0] _RAND_0;
  reg [8:0] data_reg; // @[GunzipHuffDecoder.scala 43:21:@832.4]
  reg [31:0] _RAND_1;
  wire  _T_122; // @[GunzipHuffDecoder.scala 52:19:@839.6]
  wire  _T_125; // @[GunzipHuffDecoder.scala 54:13:@842.8]
  wire [10:0] _T_128; // @[GunzipHuffDecoder.scala 58:25:@850.10]
  wire [11:0] _T_130; // @[GunzipHuffDecoder.scala 58:30:@851.10]
  wire [10:0] _T_131; // @[GunzipHuffDecoder.scala 58:30:@852.10]
  wire [10:0] _GEN_206; // @[GunzipHuffDecoder.scala 58:36:@853.10]
  wire [11:0] _T_132; // @[GunzipHuffDecoder.scala 58:36:@853.10]
  wire [10:0] _T_133; // @[GunzipHuffDecoder.scala 58:36:@854.10]
  wire [4:0] _T_135; // @[:@856.10]
  wire  _GEN_2; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire  _GEN_4; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire  _GEN_6; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire  _GEN_8; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire  _GEN_10; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire  _GEN_12; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire  _GEN_14; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire  _GEN_16; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire  _GEN_18; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire  _GEN_20; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire  _GEN_22; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire [8:0] _GEN_23; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire  _GEN_24; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire [8:0] _GEN_25; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire  _GEN_26; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire [8:0] _GEN_27; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire  _GEN_28; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire [8:0] _GEN_29; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire  _GEN_30; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire [8:0] _GEN_31; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire  _GEN_32; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire [8:0] _GEN_33; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire  _GEN_34; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire [8:0] _GEN_35; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire  _GEN_36; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire [8:0] _GEN_37; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire  _GEN_38; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire [8:0] _GEN_39; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire  _GEN_40; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire [8:0] _GEN_41; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire  _GEN_42; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire [8:0] _GEN_43; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire  _GEN_44; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire [8:0] _GEN_45; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire  _GEN_46; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire [8:0] _GEN_47; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire  _GEN_48; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire [8:0] _GEN_49; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire  _GEN_50; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire [8:0] _GEN_51; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire  _GEN_52; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire [8:0] _GEN_53; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire  _GEN_54; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire [8:0] _GEN_55; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire  _GEN_56; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire [8:0] _GEN_57; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire  _GEN_58; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire [8:0] _GEN_59; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire  _GEN_60; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire [8:0] _GEN_61; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire [10:0] _GEN_186; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire  _GEN_187; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire [8:0] _GEN_188; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  wire  _GEN_191; // @[GunzipHuffDecoder.scala 55:29:@848.8]
  wire [10:0] _GEN_192; // @[GunzipHuffDecoder.scala 55:29:@848.8]
  wire [8:0] _GEN_193; // @[GunzipHuffDecoder.scala 55:29:@848.8]
  wire  _GEN_195; // @[GunzipHuffDecoder.scala 55:29:@848.8]
  wire  _GEN_196; // @[GunzipHuffDecoder.scala 52:46:@840.6]
  wire [10:0] _GEN_197; // @[GunzipHuffDecoder.scala 52:46:@840.6]
  wire [8:0] _GEN_198; // @[GunzipHuffDecoder.scala 52:46:@840.6]
  wire  _GEN_200; // @[GunzipHuffDecoder.scala 52:46:@840.6]
  wire [10:0] _GEN_202; // @[GunzipHuffDecoder.scala 51:27:@838.4]
  wire  _GEN_207; // @[GunzipHuffDecoder.scala 54:13:@844.10]
  assign _T_122 = lit_idx >= 9'h1f; // @[GunzipHuffDecoder.scala 52:19:@839.6]
  assign _T_125 = reset == 1'h0; // @[GunzipHuffDecoder.scala 54:13:@842.8]
  assign _T_128 = lit_idx * 9'h2; // @[GunzipHuffDecoder.scala 58:25:@850.10]
  assign _T_130 = _T_128 + 11'h1; // @[GunzipHuffDecoder.scala 58:30:@851.10]
  assign _T_131 = _T_128 + 11'h1; // @[GunzipHuffDecoder.scala 58:30:@852.10]
  assign _GEN_206 = {{10'd0}, io_data_in_bits}; // @[GunzipHuffDecoder.scala 58:36:@853.10]
  assign _T_132 = _T_131 + _GEN_206; // @[GunzipHuffDecoder.scala 58:36:@853.10]
  assign _T_133 = _T_131 + _GEN_206; // @[GunzipHuffDecoder.scala 58:36:@854.10]
  assign _T_135 = lit_idx[4:0]; // @[:@856.10]
  assign _GEN_2 = 5'h1 == _T_135; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_4 = 5'h2 == _T_135 ? 1'h0 : _GEN_2; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_6 = 5'h3 == _T_135 ? 1'h0 : _GEN_4; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_8 = 5'h4 == _T_135 ? 1'h0 : _GEN_6; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_10 = 5'h5 == _T_135 ? 1'h0 : _GEN_8; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_12 = 5'h6 == _T_135 ? 1'h0 : _GEN_10; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_14 = 5'h7 == _T_135 ? 1'h0 : _GEN_12; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_16 = 5'h8 == _T_135 ? 1'h0 : _GEN_14; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_18 = 5'h9 == _T_135 ? 1'h0 : _GEN_16; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_20 = 5'ha == _T_135 ? 1'h0 : _GEN_18; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_22 = 5'hb == _T_135 ? 1'h1 : _GEN_20; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_23 = 5'hb == _T_135 ? 9'h5 : 9'h0; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_24 = 5'hc == _T_135 ? 1'h1 : _GEN_22; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_25 = 5'hc == _T_135 ? 9'h9 : _GEN_23; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_26 = 5'hd == _T_135 ? 1'h1 : _GEN_24; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_27 = 5'hd == _T_135 ? 9'he : _GEN_25; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_28 = 5'he == _T_135 ? 1'h0 : _GEN_26; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_29 = 5'he == _T_135 ? 9'h0 : _GEN_27; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_30 = 5'hf == _T_135 ? 1'h0 : _GEN_28; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_31 = 5'hf == _T_135 ? 9'h0 : _GEN_29; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_32 = 5'h10 == _T_135 ? 1'h0 : _GEN_30; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_33 = 5'h10 == _T_135 ? 9'h0 : _GEN_31; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_34 = 5'h11 == _T_135 ? 1'h0 : _GEN_32; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_35 = 5'h11 == _T_135 ? 9'h0 : _GEN_33; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_36 = 5'h12 == _T_135 ? 1'h0 : _GEN_34; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_37 = 5'h12 == _T_135 ? 9'h0 : _GEN_35; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_38 = 5'h13 == _T_135 ? 1'h0 : _GEN_36; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_39 = 5'h13 == _T_135 ? 9'h0 : _GEN_37; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_40 = 5'h14 == _T_135 ? 1'h0 : _GEN_38; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_41 = 5'h14 == _T_135 ? 9'h0 : _GEN_39; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_42 = 5'h15 == _T_135 ? 1'h0 : _GEN_40; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_43 = 5'h15 == _T_135 ? 9'h0 : _GEN_41; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_44 = 5'h16 == _T_135 ? 1'h0 : _GEN_42; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_45 = 5'h16 == _T_135 ? 9'h0 : _GEN_43; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_46 = 5'h17 == _T_135 ? 1'h0 : _GEN_44; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_47 = 5'h17 == _T_135 ? 9'h0 : _GEN_45; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_48 = 5'h18 == _T_135 ? 1'h0 : _GEN_46; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_49 = 5'h18 == _T_135 ? 9'h0 : _GEN_47; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_50 = 5'h19 == _T_135 ? 1'h0 : _GEN_48; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_51 = 5'h19 == _T_135 ? 9'h0 : _GEN_49; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_52 = 5'h1a == _T_135 ? 1'h0 : _GEN_50; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_53 = 5'h1a == _T_135 ? 9'h0 : _GEN_51; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_54 = 5'h1b == _T_135 ? 1'h0 : _GEN_52; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_55 = 5'h1b == _T_135 ? 9'h0 : _GEN_53; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_56 = 5'h1c == _T_135 ? 1'h0 : _GEN_54; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_57 = 5'h1c == _T_135 ? 9'h0 : _GEN_55; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_58 = 5'h1d == _T_135 ? 1'h1 : _GEN_56; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_59 = 5'h1d == _T_135 ? 9'h8 : _GEN_57; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_60 = 5'h1e == _T_135 ? 1'h1 : _GEN_58; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_61 = 5'h1e == _T_135 ? 9'ha : _GEN_59; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_186 = _GEN_60 ? 11'h0 : _T_133; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_187 = _GEN_60 ? 1'h0 : 1'h1; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_188 = _GEN_60 ? _GEN_61 : data_reg; // @[GunzipHuffDecoder.scala 60:43:@857.10]
  assign _GEN_191 = io_enable ? _GEN_187 : 1'h0; // @[GunzipHuffDecoder.scala 55:29:@848.8]
  assign _GEN_192 = io_enable ? _GEN_186 : 11'h0; // @[GunzipHuffDecoder.scala 55:29:@848.8]
  assign _GEN_193 = io_enable ? _GEN_188 : data_reg; // @[GunzipHuffDecoder.scala 55:29:@848.8]
  assign _GEN_195 = io_enable ? _GEN_60 : 1'h0; // @[GunzipHuffDecoder.scala 55:29:@848.8]
  assign _GEN_196 = _T_122 ? 1'h0 : _GEN_191; // @[GunzipHuffDecoder.scala 52:46:@840.6]
  assign _GEN_197 = _T_122 ? {{2'd0}, lit_idx} : _GEN_192; // @[GunzipHuffDecoder.scala 52:46:@840.6]
  assign _GEN_198 = _T_122 ? data_reg : _GEN_193; // @[GunzipHuffDecoder.scala 52:46:@840.6]
  assign _GEN_200 = _T_122 ? 1'h0 : _GEN_195; // @[GunzipHuffDecoder.scala 52:46:@840.6]
  assign _GEN_202 = io_data_in_valid ? _GEN_197 : {{2'd0}, lit_idx}; // @[GunzipHuffDecoder.scala 51:27:@838.4]
  assign io_data_in_ready = io_data_in_valid ? _GEN_196 : 1'h0; // @[GunzipHuffDecoder.scala 46:20:@835.4 GunzipHuffDecoder.scala 56:24:@849.10 GunzipHuffDecoder.scala 62:26:@859.12]
  assign io_data = io_data_in_valid ? _GEN_198 : data_reg; // @[GunzipHuffDecoder.scala 48:11:@836.4 GunzipHuffDecoder.scala 63:17:@861.12]
  assign io_valid = io_data_in_valid ? _GEN_200 : 1'h0; // @[GunzipHuffDecoder.scala 49:12:@837.4 GunzipHuffDecoder.scala 65:18:@864.12]
  assign _GEN_207 = io_data_in_valid & _T_122; // @[GunzipHuffDecoder.scala 54:13:@844.10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lit_idx = _RAND_0[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  data_reg = _RAND_1[8:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      lit_idx <= 9'h0;
    end else begin
      lit_idx <= _GEN_202[8:0];
    end
    if (io_data_in_valid) begin
      if (!(_T_122)) begin
        if (io_enable) begin
          if (_GEN_60) begin
            if (5'h1e == _T_135) begin
              data_reg <= 9'ha;
            end else begin
              if (5'h1d == _T_135) begin
                data_reg <= 9'h8;
              end else begin
                if (5'h1c == _T_135) begin
                  data_reg <= 9'h0;
                end else begin
                  if (5'h1b == _T_135) begin
                    data_reg <= 9'h0;
                  end else begin
                    if (5'h1a == _T_135) begin
                      data_reg <= 9'h0;
                    end else begin
                      if (5'h19 == _T_135) begin
                        data_reg <= 9'h0;
                      end else begin
                        if (5'h18 == _T_135) begin
                          data_reg <= 9'h0;
                        end else begin
                          if (5'h17 == _T_135) begin
                            data_reg <= 9'h0;
                          end else begin
                            if (5'h16 == _T_135) begin
                              data_reg <= 9'h0;
                            end else begin
                              if (5'h15 == _T_135) begin
                                data_reg <= 9'h0;
                              end else begin
                                if (5'h14 == _T_135) begin
                                  data_reg <= 9'h0;
                                end else begin
                                  if (5'h13 == _T_135) begin
                                    data_reg <= 9'h0;
                                  end else begin
                                    if (5'h12 == _T_135) begin
                                      data_reg <= 9'h0;
                                    end else begin
                                      if (5'h11 == _T_135) begin
                                        data_reg <= 9'h0;
                                      end else begin
                                        if (5'h10 == _T_135) begin
                                          data_reg <= 9'h0;
                                        end else begin
                                          if (5'hf == _T_135) begin
                                            data_reg <= 9'h0;
                                          end else begin
                                            if (5'he == _T_135) begin
                                              data_reg <= 9'h0;
                                            end else begin
                                              if (5'hd == _T_135) begin
                                                data_reg <= 9'he;
                                              end else begin
                                                if (5'hc == _T_135) begin
                                                  data_reg <= 9'h9;
                                                end else begin
                                                  if (5'hb == _T_135) begin
                                                    data_reg <= 9'h5;
                                                  end else begin
                                                    data_reg <= 9'h0;
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_207 & _T_125) begin
          $fwrite(32'h80000002,"DEC ERR\n"); // @[GunzipHuffDecoder.scala 54:13:@844.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module GunzipLenDistLut_1( // @[:@872.2]
  input         clock, // @[:@873.4]
  input         reset, // @[:@874.4]
  input         io_data_in_valid, // @[:@875.4]
  output        io_data_in_ready, // @[:@875.4]
  input         io_data_in_bits, // @[:@875.4]
  input         io_enable, // @[:@875.4]
  input  [8:0]  io_lut_idx, // @[:@875.4]
  output        io_done, // @[:@875.4]
  output [14:0] io_lut_out // @[:@875.4]
);
  reg [1:0] state; // @[GunzipLenDistLut.scala 66:22:@939.4]
  reg [31:0] _RAND_0;
  reg  done_reg; // @[GunzipLenDistLut.scala 69:21:@940.4]
  reg [31:0] _RAND_1;
  reg [14:0] out_reg; // @[GunzipLenDistLut.scala 70:20:@941.4]
  reg [31:0] _RAND_2;
  reg [8:0] val_init; // @[GunzipLenDistLut.scala 75:22:@944.4]
  reg [31:0] _RAND_3;
  reg [4:0] ext_idx; // @[GunzipLenDistLut.scala 76:21:@945.4]
  reg [31:0] _RAND_4;
  reg [4:0] ext_lim; // @[GunzipLenDistLut.scala 77:21:@946.4]
  reg [31:0] _RAND_5;
  reg [6:0] ext_val; // @[GunzipLenDistLut.scala 78:21:@947.4]
  reg [31:0] _RAND_6;
  wire  _T_158; // @[Conditional.scala 37:30:@948.4]
  wire  _T_160; // @[GunzipLenDistLut.scala 82:26:@950.6]
  wire  _T_161; // @[GunzipLenDistLut.scala 82:23:@951.6]
  wire [4:0] _T_163; // @[:@953.8]
  wire [14:0] _GEN_4; // @[GunzipLenDistLut.scala 83:32:@954.8]
  wire [14:0] _GEN_5; // @[GunzipLenDistLut.scala 83:32:@954.8]
  wire [14:0] _GEN_6; // @[GunzipLenDistLut.scala 83:32:@954.8]
  wire [14:0] _GEN_7; // @[GunzipLenDistLut.scala 83:32:@954.8]
  wire [14:0] _GEN_8; // @[GunzipLenDistLut.scala 83:32:@954.8]
  wire [14:0] _GEN_9; // @[GunzipLenDistLut.scala 83:32:@954.8]
  wire [14:0] _GEN_10; // @[GunzipLenDistLut.scala 83:32:@954.8]
  wire [14:0] _GEN_11; // @[GunzipLenDistLut.scala 83:32:@954.8]
  wire [14:0] _GEN_12; // @[GunzipLenDistLut.scala 83:32:@954.8]
  wire [14:0] _GEN_13; // @[GunzipLenDistLut.scala 83:32:@954.8]
  wire [14:0] _GEN_14; // @[GunzipLenDistLut.scala 83:32:@954.8]
  wire [14:0] _GEN_15; // @[GunzipLenDistLut.scala 83:32:@954.8]
  wire [14:0] _GEN_16; // @[GunzipLenDistLut.scala 83:32:@954.8]
  wire [14:0] _GEN_17; // @[GunzipLenDistLut.scala 83:32:@954.8]
  wire [14:0] _GEN_18; // @[GunzipLenDistLut.scala 83:32:@954.8]
  wire [14:0] _GEN_19; // @[GunzipLenDistLut.scala 83:32:@954.8]
  wire [14:0] _GEN_20; // @[GunzipLenDistLut.scala 83:32:@954.8]
  wire [14:0] _GEN_21; // @[GunzipLenDistLut.scala 83:32:@954.8]
  wire [14:0] _GEN_22; // @[GunzipLenDistLut.scala 83:32:@954.8]
  wire [14:0] _GEN_23; // @[GunzipLenDistLut.scala 83:32:@954.8]
  wire [14:0] _GEN_24; // @[GunzipLenDistLut.scala 83:32:@954.8]
  wire [14:0] _GEN_25; // @[GunzipLenDistLut.scala 83:32:@954.8]
  wire [14:0] _GEN_26; // @[GunzipLenDistLut.scala 83:32:@954.8]
  wire [14:0] _GEN_27; // @[GunzipLenDistLut.scala 83:32:@954.8]
  wire [14:0] _GEN_28; // @[GunzipLenDistLut.scala 83:32:@954.8]
  wire [14:0] _GEN_29; // @[GunzipLenDistLut.scala 83:32:@954.8]
  wire  _T_165; // @[GunzipLenDistLut.scala 83:32:@954.8]
  wire [14:0] _GEN_31; // @[GunzipLenDistLut.scala 85:20:@958.10]
  wire [14:0] _GEN_32; // @[GunzipLenDistLut.scala 85:20:@958.10]
  wire [14:0] _GEN_33; // @[GunzipLenDistLut.scala 85:20:@958.10]
  wire [14:0] _GEN_34; // @[GunzipLenDistLut.scala 85:20:@958.10]
  wire [14:0] _GEN_35; // @[GunzipLenDistLut.scala 85:20:@958.10]
  wire [14:0] _GEN_36; // @[GunzipLenDistLut.scala 85:20:@958.10]
  wire [14:0] _GEN_37; // @[GunzipLenDistLut.scala 85:20:@958.10]
  wire [14:0] _GEN_38; // @[GunzipLenDistLut.scala 85:20:@958.10]
  wire [14:0] _GEN_39; // @[GunzipLenDistLut.scala 85:20:@958.10]
  wire [14:0] _GEN_40; // @[GunzipLenDistLut.scala 85:20:@958.10]
  wire [14:0] _GEN_41; // @[GunzipLenDistLut.scala 85:20:@958.10]
  wire [14:0] _GEN_42; // @[GunzipLenDistLut.scala 85:20:@958.10]
  wire [14:0] _GEN_43; // @[GunzipLenDistLut.scala 85:20:@958.10]
  wire [14:0] _GEN_44; // @[GunzipLenDistLut.scala 85:20:@958.10]
  wire [14:0] _GEN_45; // @[GunzipLenDistLut.scala 85:20:@958.10]
  wire [14:0] _GEN_46; // @[GunzipLenDistLut.scala 85:20:@958.10]
  wire [14:0] _GEN_47; // @[GunzipLenDistLut.scala 85:20:@958.10]
  wire [14:0] _GEN_48; // @[GunzipLenDistLut.scala 85:20:@958.10]
  wire [14:0] _GEN_49; // @[GunzipLenDistLut.scala 85:20:@958.10]
  wire [14:0] _GEN_50; // @[GunzipLenDistLut.scala 85:20:@958.10]
  wire [14:0] _GEN_51; // @[GunzipLenDistLut.scala 85:20:@958.10]
  wire [14:0] _GEN_52; // @[GunzipLenDistLut.scala 85:20:@958.10]
  wire [14:0] _GEN_53; // @[GunzipLenDistLut.scala 85:20:@958.10]
  wire [14:0] _GEN_54; // @[GunzipLenDistLut.scala 85:20:@958.10]
  wire [14:0] _GEN_55; // @[GunzipLenDistLut.scala 85:20:@958.10]
  wire [14:0] _GEN_56; // @[GunzipLenDistLut.scala 85:20:@958.10]
  wire [14:0] _GEN_57; // @[GunzipLenDistLut.scala 85:20:@958.10]
  wire [14:0] _GEN_58; // @[GunzipLenDistLut.scala 85:20:@958.10]
  wire [14:0] _GEN_59; // @[GunzipLenDistLut.scala 85:20:@958.10]
  wire [15:0] _T_172; // @[GunzipLenDistLut.scala 87:39:@961.10]
  wire [15:0] _T_173; // @[GunzipLenDistLut.scala 87:39:@962.10]
  wire [14:0] _T_174; // @[GunzipLenDistLut.scala 87:39:@963.10]
  wire [1:0] _GEN_120; // @[GunzipLenDistLut.scala 83:39:@955.8]
  wire [14:0] _GEN_121; // @[GunzipLenDistLut.scala 83:39:@955.8]
  wire [4:0] _GEN_122; // @[GunzipLenDistLut.scala 83:39:@955.8]
  wire [14:0] _GEN_123; // @[GunzipLenDistLut.scala 83:39:@955.8]
  wire [6:0] _GEN_124; // @[GunzipLenDistLut.scala 83:39:@955.8]
  wire  _GEN_125; // @[GunzipLenDistLut.scala 83:39:@955.8]
  wire [14:0] _GEN_126; // @[GunzipLenDistLut.scala 83:39:@955.8]
  wire [1:0] _GEN_127; // @[GunzipLenDistLut.scala 82:36:@952.6]
  wire [14:0] _GEN_128; // @[GunzipLenDistLut.scala 82:36:@952.6]
  wire [4:0] _GEN_129; // @[GunzipLenDistLut.scala 82:36:@952.6]
  wire [14:0] _GEN_130; // @[GunzipLenDistLut.scala 82:36:@952.6]
  wire [6:0] _GEN_131; // @[GunzipLenDistLut.scala 82:36:@952.6]
  wire  _GEN_132; // @[GunzipLenDistLut.scala 82:36:@952.6]
  wire [14:0] _GEN_133; // @[GunzipLenDistLut.scala 82:36:@952.6]
  wire  _T_179; // @[Conditional.scala 37:30:@976.6]
  wire  _T_185; // @[Conditional.scala 37:30:@982.10]
  wire [5:0] _T_186; // @[GunzipLenDistLut.scala 50:33:@984.12]
  wire [6:0] _T_187; // @[Cat.scala 30:58:@985.12]
  wire  _T_189; // @[Conditional.scala 37:30:@989.12]
  wire [4:0] _T_190; // @[GunzipLenDistLut.scala 51:33:@991.14]
  wire  _T_191; // @[GunzipLenDistLut.scala 51:70:@992.14]
  wire [6:0] _T_193; // @[Cat.scala 30:58:@994.14]
  wire  _T_195; // @[Conditional.scala 37:30:@998.14]
  wire [3:0] _T_196; // @[GunzipLenDistLut.scala 52:33:@1000.16]
  wire [1:0] _T_197; // @[GunzipLenDistLut.scala 52:70:@1001.16]
  wire [6:0] _T_199; // @[Cat.scala 30:58:@1003.16]
  wire  _T_201; // @[Conditional.scala 37:30:@1007.16]
  wire [2:0] _T_202; // @[GunzipLenDistLut.scala 53:33:@1009.18]
  wire [2:0] _T_203; // @[GunzipLenDistLut.scala 53:70:@1010.18]
  wire [6:0] _T_205; // @[Cat.scala 30:58:@1012.18]
  wire  _T_207; // @[Conditional.scala 37:30:@1016.18]
  wire [1:0] _T_208; // @[GunzipLenDistLut.scala 54:33:@1018.20]
  wire [3:0] _T_209; // @[GunzipLenDistLut.scala 54:70:@1019.20]
  wire [6:0] _T_211; // @[Cat.scala 30:58:@1021.20]
  wire  _T_213; // @[Conditional.scala 37:30:@1025.20]
  wire  _T_214; // @[GunzipLenDistLut.scala 55:33:@1027.22]
  wire [4:0] _T_215; // @[GunzipLenDistLut.scala 55:70:@1028.22]
  wire [6:0] _T_217; // @[Cat.scala 30:58:@1030.22]
  wire [6:0] _GEN_134; // @[Conditional.scala 39:67:@1026.20]
  wire [6:0] _GEN_135; // @[Conditional.scala 39:67:@1017.18]
  wire [6:0] _GEN_136; // @[Conditional.scala 39:67:@1008.16]
  wire [6:0] _GEN_137; // @[Conditional.scala 39:67:@999.14]
  wire [6:0] _GEN_138; // @[Conditional.scala 39:67:@990.12]
  wire [6:0] _GEN_139; // @[Conditional.scala 40:58:@983.10]
  wire [5:0] _T_219; // @[GunzipLenDistLut.scala 100:28:@1034.10]
  wire [4:0] _T_220; // @[GunzipLenDistLut.scala 100:28:@1035.10]
  wire  _T_221; // @[GunzipLenDistLut.scala 102:22:@1037.10]
  wire [1:0] _GEN_140; // @[GunzipLenDistLut.scala 102:35:@1038.10]
  wire [6:0] _GEN_142; // @[GunzipLenDistLut.scala 97:31:@978.8]
  wire [4:0] _GEN_143; // @[GunzipLenDistLut.scala 97:31:@978.8]
  wire [1:0] _GEN_144; // @[GunzipLenDistLut.scala 97:31:@978.8]
  wire  _T_222; // @[Conditional.scala 37:30:@1044.8]
  wire [8:0] _GEN_163; // @[GunzipLenDistLut.scala 110:27:@1048.10]
  wire [9:0] _T_224; // @[GunzipLenDistLut.scala 110:27:@1048.10]
  wire [8:0] _T_225; // @[GunzipLenDistLut.scala 110:27:@1049.10]
  wire [1:0] _GEN_145; // @[Conditional.scala 39:67:@1045.8]
  wire [14:0] _GEN_147; // @[Conditional.scala 39:67:@1045.8]
  wire  _GEN_148; // @[Conditional.scala 39:67:@977.6]
  wire [6:0] _GEN_149; // @[Conditional.scala 39:67:@977.6]
  wire [4:0] _GEN_150; // @[Conditional.scala 39:67:@977.6]
  wire [1:0] _GEN_151; // @[Conditional.scala 39:67:@977.6]
  wire  _GEN_152; // @[Conditional.scala 39:67:@977.6]
  wire [14:0] _GEN_153; // @[Conditional.scala 39:67:@977.6]
  wire [1:0] _GEN_154; // @[Conditional.scala 40:58:@949.4]
  wire [14:0] _GEN_155; // @[Conditional.scala 40:58:@949.4]
  wire [14:0] _GEN_157; // @[Conditional.scala 40:58:@949.4]
  wire  _GEN_161; // @[Conditional.scala 40:58:@949.4]
  assign _T_158 = 2'h0 == state; // @[Conditional.scala 37:30:@948.4]
  assign _T_160 = io_done == 1'h0; // @[GunzipLenDistLut.scala 82:26:@950.6]
  assign _T_161 = io_enable & _T_160; // @[GunzipLenDistLut.scala 82:23:@951.6]
  assign _T_163 = io_lut_idx[4:0]; // @[:@953.8]
  assign _GEN_4 = 5'h4 == _T_163 ? 15'h1 : 15'h0; // @[GunzipLenDistLut.scala 83:32:@954.8]
  assign _GEN_5 = 5'h5 == _T_163 ? 15'h1 : _GEN_4; // @[GunzipLenDistLut.scala 83:32:@954.8]
  assign _GEN_6 = 5'h6 == _T_163 ? 15'h2 : _GEN_5; // @[GunzipLenDistLut.scala 83:32:@954.8]
  assign _GEN_7 = 5'h7 == _T_163 ? 15'h2 : _GEN_6; // @[GunzipLenDistLut.scala 83:32:@954.8]
  assign _GEN_8 = 5'h8 == _T_163 ? 15'h3 : _GEN_7; // @[GunzipLenDistLut.scala 83:32:@954.8]
  assign _GEN_9 = 5'h9 == _T_163 ? 15'h3 : _GEN_8; // @[GunzipLenDistLut.scala 83:32:@954.8]
  assign _GEN_10 = 5'ha == _T_163 ? 15'h4 : _GEN_9; // @[GunzipLenDistLut.scala 83:32:@954.8]
  assign _GEN_11 = 5'hb == _T_163 ? 15'h4 : _GEN_10; // @[GunzipLenDistLut.scala 83:32:@954.8]
  assign _GEN_12 = 5'hc == _T_163 ? 15'h5 : _GEN_11; // @[GunzipLenDistLut.scala 83:32:@954.8]
  assign _GEN_13 = 5'hd == _T_163 ? 15'h5 : _GEN_12; // @[GunzipLenDistLut.scala 83:32:@954.8]
  assign _GEN_14 = 5'he == _T_163 ? 15'h6 : _GEN_13; // @[GunzipLenDistLut.scala 83:32:@954.8]
  assign _GEN_15 = 5'hf == _T_163 ? 15'h6 : _GEN_14; // @[GunzipLenDistLut.scala 83:32:@954.8]
  assign _GEN_16 = 5'h10 == _T_163 ? 15'h7 : _GEN_15; // @[GunzipLenDistLut.scala 83:32:@954.8]
  assign _GEN_17 = 5'h11 == _T_163 ? 15'h7 : _GEN_16; // @[GunzipLenDistLut.scala 83:32:@954.8]
  assign _GEN_18 = 5'h12 == _T_163 ? 15'h8 : _GEN_17; // @[GunzipLenDistLut.scala 83:32:@954.8]
  assign _GEN_19 = 5'h13 == _T_163 ? 15'h8 : _GEN_18; // @[GunzipLenDistLut.scala 83:32:@954.8]
  assign _GEN_20 = 5'h14 == _T_163 ? 15'h9 : _GEN_19; // @[GunzipLenDistLut.scala 83:32:@954.8]
  assign _GEN_21 = 5'h15 == _T_163 ? 15'h9 : _GEN_20; // @[GunzipLenDistLut.scala 83:32:@954.8]
  assign _GEN_22 = 5'h16 == _T_163 ? 15'ha : _GEN_21; // @[GunzipLenDistLut.scala 83:32:@954.8]
  assign _GEN_23 = 5'h17 == _T_163 ? 15'ha : _GEN_22; // @[GunzipLenDistLut.scala 83:32:@954.8]
  assign _GEN_24 = 5'h18 == _T_163 ? 15'hb : _GEN_23; // @[GunzipLenDistLut.scala 83:32:@954.8]
  assign _GEN_25 = 5'h19 == _T_163 ? 15'hb : _GEN_24; // @[GunzipLenDistLut.scala 83:32:@954.8]
  assign _GEN_26 = 5'h1a == _T_163 ? 15'hc : _GEN_25; // @[GunzipLenDistLut.scala 83:32:@954.8]
  assign _GEN_27 = 5'h1b == _T_163 ? 15'hc : _GEN_26; // @[GunzipLenDistLut.scala 83:32:@954.8]
  assign _GEN_28 = 5'h1c == _T_163 ? 15'hd : _GEN_27; // @[GunzipLenDistLut.scala 83:32:@954.8]
  assign _GEN_29 = 5'h1d == _T_163 ? 15'hd : _GEN_28; // @[GunzipLenDistLut.scala 83:32:@954.8]
  assign _T_165 = _GEN_29 > 15'h0; // @[GunzipLenDistLut.scala 83:32:@954.8]
  assign _GEN_31 = 5'h1 == _T_163 ? 15'h2 : 15'h1; // @[GunzipLenDistLut.scala 85:20:@958.10]
  assign _GEN_32 = 5'h2 == _T_163 ? 15'h3 : _GEN_31; // @[GunzipLenDistLut.scala 85:20:@958.10]
  assign _GEN_33 = 5'h3 == _T_163 ? 15'h4 : _GEN_32; // @[GunzipLenDistLut.scala 85:20:@958.10]
  assign _GEN_34 = 5'h4 == _T_163 ? 15'h5 : _GEN_33; // @[GunzipLenDistLut.scala 85:20:@958.10]
  assign _GEN_35 = 5'h5 == _T_163 ? 15'h7 : _GEN_34; // @[GunzipLenDistLut.scala 85:20:@958.10]
  assign _GEN_36 = 5'h6 == _T_163 ? 15'h9 : _GEN_35; // @[GunzipLenDistLut.scala 85:20:@958.10]
  assign _GEN_37 = 5'h7 == _T_163 ? 15'hd : _GEN_36; // @[GunzipLenDistLut.scala 85:20:@958.10]
  assign _GEN_38 = 5'h8 == _T_163 ? 15'h11 : _GEN_37; // @[GunzipLenDistLut.scala 85:20:@958.10]
  assign _GEN_39 = 5'h9 == _T_163 ? 15'h19 : _GEN_38; // @[GunzipLenDistLut.scala 85:20:@958.10]
  assign _GEN_40 = 5'ha == _T_163 ? 15'h21 : _GEN_39; // @[GunzipLenDistLut.scala 85:20:@958.10]
  assign _GEN_41 = 5'hb == _T_163 ? 15'h31 : _GEN_40; // @[GunzipLenDistLut.scala 85:20:@958.10]
  assign _GEN_42 = 5'hc == _T_163 ? 15'h41 : _GEN_41; // @[GunzipLenDistLut.scala 85:20:@958.10]
  assign _GEN_43 = 5'hd == _T_163 ? 15'h61 : _GEN_42; // @[GunzipLenDistLut.scala 85:20:@958.10]
  assign _GEN_44 = 5'he == _T_163 ? 15'h81 : _GEN_43; // @[GunzipLenDistLut.scala 85:20:@958.10]
  assign _GEN_45 = 5'hf == _T_163 ? 15'hc1 : _GEN_44; // @[GunzipLenDistLut.scala 85:20:@958.10]
  assign _GEN_46 = 5'h10 == _T_163 ? 15'h101 : _GEN_45; // @[GunzipLenDistLut.scala 85:20:@958.10]
  assign _GEN_47 = 5'h11 == _T_163 ? 15'h181 : _GEN_46; // @[GunzipLenDistLut.scala 85:20:@958.10]
  assign _GEN_48 = 5'h12 == _T_163 ? 15'h201 : _GEN_47; // @[GunzipLenDistLut.scala 85:20:@958.10]
  assign _GEN_49 = 5'h13 == _T_163 ? 15'h301 : _GEN_48; // @[GunzipLenDistLut.scala 85:20:@958.10]
  assign _GEN_50 = 5'h14 == _T_163 ? 15'h401 : _GEN_49; // @[GunzipLenDistLut.scala 85:20:@958.10]
  assign _GEN_51 = 5'h15 == _T_163 ? 15'h601 : _GEN_50; // @[GunzipLenDistLut.scala 85:20:@958.10]
  assign _GEN_52 = 5'h16 == _T_163 ? 15'h801 : _GEN_51; // @[GunzipLenDistLut.scala 85:20:@958.10]
  assign _GEN_53 = 5'h17 == _T_163 ? 15'hc01 : _GEN_52; // @[GunzipLenDistLut.scala 85:20:@958.10]
  assign _GEN_54 = 5'h18 == _T_163 ? 15'h1001 : _GEN_53; // @[GunzipLenDistLut.scala 85:20:@958.10]
  assign _GEN_55 = 5'h19 == _T_163 ? 15'h1801 : _GEN_54; // @[GunzipLenDistLut.scala 85:20:@958.10]
  assign _GEN_56 = 5'h1a == _T_163 ? 15'h2001 : _GEN_55; // @[GunzipLenDistLut.scala 85:20:@958.10]
  assign _GEN_57 = 5'h1b == _T_163 ? 15'h3001 : _GEN_56; // @[GunzipLenDistLut.scala 85:20:@958.10]
  assign _GEN_58 = 5'h1c == _T_163 ? 15'h4001 : _GEN_57; // @[GunzipLenDistLut.scala 85:20:@958.10]
  assign _GEN_59 = 5'h1d == _T_163 ? 15'h6001 : _GEN_58; // @[GunzipLenDistLut.scala 85:20:@958.10]
  assign _T_172 = _GEN_29 - 15'h1; // @[GunzipLenDistLut.scala 87:39:@961.10]
  assign _T_173 = $unsigned(_T_172); // @[GunzipLenDistLut.scala 87:39:@962.10]
  assign _T_174 = _T_173[14:0]; // @[GunzipLenDistLut.scala 87:39:@963.10]
  assign _GEN_120 = _T_165 ? 2'h1 : 2'h0; // @[GunzipLenDistLut.scala 83:39:@955.8]
  assign _GEN_121 = _T_165 ? _GEN_59 : {{6'd0}, val_init}; // @[GunzipLenDistLut.scala 83:39:@955.8]
  assign _GEN_122 = _T_165 ? 5'h0 : ext_idx; // @[GunzipLenDistLut.scala 83:39:@955.8]
  assign _GEN_123 = _T_165 ? _T_174 : {{10'd0}, ext_lim}; // @[GunzipLenDistLut.scala 83:39:@955.8]
  assign _GEN_124 = _T_165 ? 7'h0 : ext_val; // @[GunzipLenDistLut.scala 83:39:@955.8]
  assign _GEN_125 = _T_165 ? 1'h0 : 1'h1; // @[GunzipLenDistLut.scala 83:39:@955.8]
  assign _GEN_126 = _T_165 ? out_reg : _GEN_59; // @[GunzipLenDistLut.scala 83:39:@955.8]
  assign _GEN_127 = _T_161 ? _GEN_120 : state; // @[GunzipLenDistLut.scala 82:36:@952.6]
  assign _GEN_128 = _T_161 ? _GEN_121 : {{6'd0}, val_init}; // @[GunzipLenDistLut.scala 82:36:@952.6]
  assign _GEN_129 = _T_161 ? _GEN_122 : ext_idx; // @[GunzipLenDistLut.scala 82:36:@952.6]
  assign _GEN_130 = _T_161 ? _GEN_123 : {{10'd0}, ext_lim}; // @[GunzipLenDistLut.scala 82:36:@952.6]
  assign _GEN_131 = _T_161 ? _GEN_124 : ext_val; // @[GunzipLenDistLut.scala 82:36:@952.6]
  assign _GEN_132 = _T_161 ? _GEN_125 : 1'h0; // @[GunzipLenDistLut.scala 82:36:@952.6]
  assign _GEN_133 = _T_161 ? _GEN_126 : out_reg; // @[GunzipLenDistLut.scala 82:36:@952.6]
  assign _T_179 = 2'h1 == state; // @[Conditional.scala 37:30:@976.6]
  assign _T_185 = 5'h0 == ext_idx; // @[Conditional.scala 37:30:@982.10]
  assign _T_186 = ext_val[6:1]; // @[GunzipLenDistLut.scala 50:33:@984.12]
  assign _T_187 = {_T_186,io_data_in_bits}; // @[Cat.scala 30:58:@985.12]
  assign _T_189 = 5'h1 == ext_idx; // @[Conditional.scala 37:30:@989.12]
  assign _T_190 = ext_val[6:2]; // @[GunzipLenDistLut.scala 51:33:@991.14]
  assign _T_191 = ext_val[0]; // @[GunzipLenDistLut.scala 51:70:@992.14]
  assign _T_193 = {_T_190,io_data_in_bits,_T_191}; // @[Cat.scala 30:58:@994.14]
  assign _T_195 = 5'h2 == ext_idx; // @[Conditional.scala 37:30:@998.14]
  assign _T_196 = ext_val[6:3]; // @[GunzipLenDistLut.scala 52:33:@1000.16]
  assign _T_197 = ext_val[1:0]; // @[GunzipLenDistLut.scala 52:70:@1001.16]
  assign _T_199 = {_T_196,io_data_in_bits,_T_197}; // @[Cat.scala 30:58:@1003.16]
  assign _T_201 = 5'h3 == ext_idx; // @[Conditional.scala 37:30:@1007.16]
  assign _T_202 = ext_val[6:4]; // @[GunzipLenDistLut.scala 53:33:@1009.18]
  assign _T_203 = ext_val[2:0]; // @[GunzipLenDistLut.scala 53:70:@1010.18]
  assign _T_205 = {_T_202,io_data_in_bits,_T_203}; // @[Cat.scala 30:58:@1012.18]
  assign _T_207 = 5'h4 == ext_idx; // @[Conditional.scala 37:30:@1016.18]
  assign _T_208 = ext_val[6:5]; // @[GunzipLenDistLut.scala 54:33:@1018.20]
  assign _T_209 = ext_val[3:0]; // @[GunzipLenDistLut.scala 54:70:@1019.20]
  assign _T_211 = {_T_208,io_data_in_bits,_T_209}; // @[Cat.scala 30:58:@1021.20]
  assign _T_213 = 5'h5 == ext_idx; // @[Conditional.scala 37:30:@1025.20]
  assign _T_214 = ext_val[6]; // @[GunzipLenDistLut.scala 55:33:@1027.22]
  assign _T_215 = ext_val[4:0]; // @[GunzipLenDistLut.scala 55:70:@1028.22]
  assign _T_217 = {_T_214,io_data_in_bits,_T_215}; // @[Cat.scala 30:58:@1030.22]
  assign _GEN_134 = _T_213 ? _T_217 : 7'h0; // @[Conditional.scala 39:67:@1026.20]
  assign _GEN_135 = _T_207 ? _T_211 : _GEN_134; // @[Conditional.scala 39:67:@1017.18]
  assign _GEN_136 = _T_201 ? _T_205 : _GEN_135; // @[Conditional.scala 39:67:@1008.16]
  assign _GEN_137 = _T_195 ? _T_199 : _GEN_136; // @[Conditional.scala 39:67:@999.14]
  assign _GEN_138 = _T_189 ? _T_193 : _GEN_137; // @[Conditional.scala 39:67:@990.12]
  assign _GEN_139 = _T_185 ? _T_187 : _GEN_138; // @[Conditional.scala 40:58:@983.10]
  assign _T_219 = ext_idx + 5'h1; // @[GunzipLenDistLut.scala 100:28:@1034.10]
  assign _T_220 = ext_idx + 5'h1; // @[GunzipLenDistLut.scala 100:28:@1035.10]
  assign _T_221 = ext_idx == ext_lim; // @[GunzipLenDistLut.scala 102:22:@1037.10]
  assign _GEN_140 = _T_221 ? 2'h2 : state; // @[GunzipLenDistLut.scala 102:35:@1038.10]
  assign _GEN_142 = io_data_in_valid ? _GEN_139 : ext_val; // @[GunzipLenDistLut.scala 97:31:@978.8]
  assign _GEN_143 = io_data_in_valid ? _T_220 : ext_idx; // @[GunzipLenDistLut.scala 97:31:@978.8]
  assign _GEN_144 = io_data_in_valid ? _GEN_140 : state; // @[GunzipLenDistLut.scala 97:31:@978.8]
  assign _T_222 = 2'h2 == state; // @[Conditional.scala 37:30:@1044.8]
  assign _GEN_163 = {{2'd0}, ext_val}; // @[GunzipLenDistLut.scala 110:27:@1048.10]
  assign _T_224 = val_init + _GEN_163; // @[GunzipLenDistLut.scala 110:27:@1048.10]
  assign _T_225 = val_init + _GEN_163; // @[GunzipLenDistLut.scala 110:27:@1049.10]
  assign _GEN_145 = _T_222 ? 2'h0 : state; // @[Conditional.scala 39:67:@1045.8]
  assign _GEN_147 = _T_222 ? {{6'd0}, _T_225} : out_reg; // @[Conditional.scala 39:67:@1045.8]
  assign _GEN_148 = _T_179 ? io_data_in_valid : 1'h0; // @[Conditional.scala 39:67:@977.6]
  assign _GEN_149 = _T_179 ? _GEN_142 : ext_val; // @[Conditional.scala 39:67:@977.6]
  assign _GEN_150 = _T_179 ? _GEN_143 : ext_idx; // @[Conditional.scala 39:67:@977.6]
  assign _GEN_151 = _T_179 ? _GEN_144 : _GEN_145; // @[Conditional.scala 39:67:@977.6]
  assign _GEN_152 = _T_179 ? 1'h0 : _T_222; // @[Conditional.scala 39:67:@977.6]
  assign _GEN_153 = _T_179 ? out_reg : _GEN_147; // @[Conditional.scala 39:67:@977.6]
  assign _GEN_154 = _T_158 ? _GEN_127 : _GEN_151; // @[Conditional.scala 40:58:@949.4]
  assign _GEN_155 = _T_158 ? _GEN_128 : {{6'd0}, val_init}; // @[Conditional.scala 40:58:@949.4]
  assign _GEN_157 = _T_158 ? _GEN_130 : {{10'd0}, ext_lim}; // @[Conditional.scala 40:58:@949.4]
  assign _GEN_161 = _T_158 ? 1'h0 : _GEN_148; // @[Conditional.scala 40:58:@949.4]
  assign io_data_in_ready = done_reg ? 1'h0 : _GEN_161; // @[GunzipLenDistLut.scala 72:20:@943.4 GunzipLenDistLut.scala 98:26:@979.10 GunzipLenDistLut.scala 118:22:@1055.6]
  assign io_done = done_reg; // @[GunzipLenDistLut.scala 115:11:@1053.4]
  assign io_lut_out = out_reg; // @[GunzipLenDistLut.scala 114:14:@1052.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  done_reg = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_reg = _RAND_2[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  val_init = _RAND_3[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  ext_idx = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  ext_lim = _RAND_5[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  ext_val = _RAND_6[6:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_158) begin
        if (_T_161) begin
          if (_T_165) begin
            state <= 2'h1;
          end else begin
            state <= 2'h0;
          end
        end
      end else begin
        if (_T_179) begin
          if (io_data_in_valid) begin
            if (_T_221) begin
              state <= 2'h2;
            end
          end
        end else begin
          if (_T_222) begin
            state <= 2'h0;
          end
        end
      end
    end
    if (_T_158) begin
      if (_T_161) begin
        if (_T_165) begin
          done_reg <= 1'h0;
        end else begin
          done_reg <= 1'h1;
        end
      end else begin
        done_reg <= 1'h0;
      end
    end else begin
      if (_T_179) begin
        done_reg <= 1'h0;
      end else begin
        done_reg <= _T_222;
      end
    end
    if (_T_158) begin
      if (_T_161) begin
        if (!(_T_165)) begin
          if (5'h1d == _T_163) begin
            out_reg <= 15'h6001;
          end else begin
            if (5'h1c == _T_163) begin
              out_reg <= 15'h4001;
            end else begin
              if (5'h1b == _T_163) begin
                out_reg <= 15'h3001;
              end else begin
                if (5'h1a == _T_163) begin
                  out_reg <= 15'h2001;
                end else begin
                  if (5'h19 == _T_163) begin
                    out_reg <= 15'h1801;
                  end else begin
                    if (5'h18 == _T_163) begin
                      out_reg <= 15'h1001;
                    end else begin
                      if (5'h17 == _T_163) begin
                        out_reg <= 15'hc01;
                      end else begin
                        if (5'h16 == _T_163) begin
                          out_reg <= 15'h801;
                        end else begin
                          if (5'h15 == _T_163) begin
                            out_reg <= 15'h601;
                          end else begin
                            if (5'h14 == _T_163) begin
                              out_reg <= 15'h401;
                            end else begin
                              if (5'h13 == _T_163) begin
                                out_reg <= 15'h301;
                              end else begin
                                if (5'h12 == _T_163) begin
                                  out_reg <= 15'h201;
                                end else begin
                                  if (5'h11 == _T_163) begin
                                    out_reg <= 15'h181;
                                  end else begin
                                    if (5'h10 == _T_163) begin
                                      out_reg <= 15'h101;
                                    end else begin
                                      if (5'hf == _T_163) begin
                                        out_reg <= 15'hc1;
                                      end else begin
                                        if (5'he == _T_163) begin
                                          out_reg <= 15'h81;
                                        end else begin
                                          if (5'hd == _T_163) begin
                                            out_reg <= 15'h61;
                                          end else begin
                                            if (5'hc == _T_163) begin
                                              out_reg <= 15'h41;
                                            end else begin
                                              if (5'hb == _T_163) begin
                                                out_reg <= 15'h31;
                                              end else begin
                                                if (5'ha == _T_163) begin
                                                  out_reg <= 15'h21;
                                                end else begin
                                                  if (5'h9 == _T_163) begin
                                                    out_reg <= 15'h19;
                                                  end else begin
                                                    if (5'h8 == _T_163) begin
                                                      out_reg <= 15'h11;
                                                    end else begin
                                                      if (5'h7 == _T_163) begin
                                                        out_reg <= 15'hd;
                                                      end else begin
                                                        if (5'h6 == _T_163) begin
                                                          out_reg <= 15'h9;
                                                        end else begin
                                                          if (5'h5 == _T_163) begin
                                                            out_reg <= 15'h7;
                                                          end else begin
                                                            if (5'h4 == _T_163) begin
                                                              out_reg <= 15'h5;
                                                            end else begin
                                                              if (5'h3 == _T_163) begin
                                                                out_reg <= 15'h4;
                                                              end else begin
                                                                if (5'h2 == _T_163) begin
                                                                  out_reg <= 15'h3;
                                                                end else begin
                                                                  if (5'h1 == _T_163) begin
                                                                    out_reg <= 15'h2;
                                                                  end else begin
                                                                    out_reg <= 15'h1;
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (!(_T_179)) begin
        if (_T_222) begin
          out_reg <= {{6'd0}, _T_225};
        end
      end
    end
    val_init <= _GEN_155[8:0];
    if (_T_158) begin
      if (_T_161) begin
        if (_T_165) begin
          ext_idx <= 5'h0;
        end
      end
    end else begin
      if (_T_179) begin
        if (io_data_in_valid) begin
          ext_idx <= _T_220;
        end
      end
    end
    ext_lim <= _GEN_157[4:0];
    if (_T_158) begin
      if (_T_161) begin
        if (_T_165) begin
          ext_val <= 7'h0;
        end
      end
    end else begin
      if (_T_179) begin
        if (io_data_in_valid) begin
          if (_T_185) begin
            ext_val <= _T_187;
          end else begin
            if (_T_189) begin
              ext_val <= _T_193;
            end else begin
              if (_T_195) begin
                ext_val <= _T_199;
              end else begin
                if (_T_201) begin
                  ext_val <= _T_205;
                end else begin
                  if (_T_207) begin
                    ext_val <= _T_211;
                  end else begin
                    if (_T_213) begin
                      ext_val <= _T_217;
                    end else begin
                      ext_val <= 7'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
  end
endmodule
module GunzipOutBuf( // @[:@1058.2]
  input         clock, // @[:@1059.4]
  input         reset, // @[:@1060.4]
  input  [7:0]  io_data_in, // @[:@1061.4]
  input         io_valid_in, // @[:@1061.4]
  input  [14:0] io_dist, // @[:@1061.4]
  input  [14:0] io_len, // @[:@1061.4]
  input         io_enable, // @[:@1061.4]
  output        io_done, // @[:@1061.4]
  output [7:0]  io_data_out_bits, // @[:@1061.4]
  output        io_data_out_valid, // @[:@1061.4]
  input         io_data_out_ready // @[:@1061.4]
);
  reg [7:0] out_buf [0:32767]; // @[GunzipOutBuf.scala 46:28:@1063.4]
  reg [31:0] _RAND_0;
  wire [7:0] out_buf__T_59_data; // @[GunzipOutBuf.scala 46:28:@1063.4]
  wire [14:0] out_buf__T_59_addr; // @[GunzipOutBuf.scala 46:28:@1063.4]
  wire [7:0] out_buf__T_30_data; // @[GunzipOutBuf.scala 46:28:@1063.4]
  wire [14:0] out_buf__T_30_addr; // @[GunzipOutBuf.scala 46:28:@1063.4]
  wire  out_buf__T_30_mask; // @[GunzipOutBuf.scala 46:28:@1063.4]
  wire  out_buf__T_30_en; // @[GunzipOutBuf.scala 46:28:@1063.4]
  reg [14:0] out_buf_wr_pos; // @[GunzipOutBuf.scala 47:31:@1064.4]
  reg [31:0] _RAND_1;
  reg [14:0] out_buf_rd_pos; // @[GunzipOutBuf.scala 48:31:@1065.4]
  reg [31:0] _RAND_2;
  reg [14:0] rem_len; // @[GunzipOutBuf.scala 49:20:@1066.4]
  reg [31:0] _RAND_3;
  wire [15:0] _T_32; // @[GunzipOutBuf.scala 54:38:@1070.6]
  wire [14:0] _T_33; // @[GunzipOutBuf.scala 54:38:@1071.6]
  wire  _GEN_3; // @[GunzipOutBuf.scala 52:22:@1067.4]
  wire [14:0] _GEN_5; // @[GunzipOutBuf.scala 52:22:@1067.4]
  reg [1:0] state; // @[GunzipOutBuf.scala 58:22:@1074.4]
  reg [31:0] _RAND_4;
  wire  _T_35; // @[Conditional.scala 37:30:@1075.4]
  wire [1:0] _GEN_6; // @[GunzipOutBuf.scala 62:24:@1077.6]
  wire  _T_36; // @[Conditional.scala 37:30:@1082.6]
  wire  _T_37; // @[Conditional.scala 37:30:@1087.8]
  wire [1:0] _GEN_7; // @[GunzipOutBuf.scala 70:32:@1089.10]
  wire  _T_38; // @[Conditional.scala 37:30:@1094.10]
  wire [1:0] _GEN_8; // @[GunzipOutBuf.scala 75:22:@1096.12]
  wire [1:0] _GEN_9; // @[Conditional.scala 39:67:@1095.10]
  wire [1:0] _GEN_10; // @[Conditional.scala 39:67:@1088.8]
  wire [1:0] _GEN_11; // @[Conditional.scala 39:67:@1083.6]
  wire [1:0] _GEN_12; // @[Conditional.scala 40:58:@1076.4]
  wire  _T_39; // @[GunzipOutBuf.scala 83:15:@1103.4]
  wire  _T_40; // @[GunzipOutBuf.scala 83:25:@1104.4]
  wire [15:0] _T_41; // @[GunzipOutBuf.scala 84:38:@1106.6]
  wire [15:0] _T_42; // @[GunzipOutBuf.scala 84:38:@1107.6]
  wire [14:0] _T_43; // @[GunzipOutBuf.scala 84:38:@1108.6]
  wire  _T_44; // @[GunzipOutBuf.scala 86:22:@1113.6]
  wire  _T_45; // @[GunzipOutBuf.scala 86:32:@1114.6]
  wire [15:0] _T_47; // @[GunzipOutBuf.scala 87:38:@1116.8]
  wire [14:0] _T_48; // @[GunzipOutBuf.scala 87:38:@1117.8]
  wire [15:0] _T_50; // @[GunzipOutBuf.scala 88:24:@1119.8]
  wire [15:0] _T_51; // @[GunzipOutBuf.scala 88:24:@1120.8]
  wire [14:0] _T_52; // @[GunzipOutBuf.scala 88:24:@1121.8]
  wire [14:0] _GEN_13; // @[GunzipOutBuf.scala 86:54:@1115.6]
  wire [14:0] _GEN_14; // @[GunzipOutBuf.scala 86:54:@1115.6]
  wire [14:0] _GEN_15; // @[GunzipOutBuf.scala 83:39:@1105.4]
  wire  _T_61; // @[GunzipOutBuf.scala 94:20:@1135.4]
  wire  _T_63; // @[GunzipOutBuf.scala 94:42:@1136.4]
  reg [14:0] out_buf__T_59_addr_pipe_0;
  reg [31:0] _RAND_5;
  assign out_buf__T_59_addr = out_buf__T_59_addr_pipe_0;
  assign out_buf__T_59_data = out_buf[out_buf__T_59_addr]; // @[GunzipOutBuf.scala 46:28:@1063.4]
  assign out_buf__T_30_data = io_data_in;
  assign out_buf__T_30_addr = out_buf_wr_pos;
  assign out_buf__T_30_mask = 1'h1;
  assign out_buf__T_30_en = io_valid_in;
  assign _T_32 = out_buf_wr_pos + 15'h1; // @[GunzipOutBuf.scala 54:38:@1070.6]
  assign _T_33 = out_buf_wr_pos + 15'h1; // @[GunzipOutBuf.scala 54:38:@1071.6]
  assign _GEN_3 = 1'h1; // @[GunzipOutBuf.scala 52:22:@1067.4]
  assign _GEN_5 = io_valid_in ? _T_33 : out_buf_wr_pos; // @[GunzipOutBuf.scala 52:22:@1067.4]
  assign _T_35 = 2'h0 == state; // @[Conditional.scala 37:30:@1075.4]
  assign _GEN_6 = io_enable ? 2'h1 : state; // @[GunzipOutBuf.scala 62:24:@1077.6]
  assign _T_36 = 2'h1 == state; // @[Conditional.scala 37:30:@1082.6]
  assign _T_37 = 2'h2 == state; // @[Conditional.scala 37:30:@1087.8]
  assign _GEN_7 = io_data_out_ready ? 2'h3 : state; // @[GunzipOutBuf.scala 70:32:@1089.10]
  assign _T_38 = 2'h3 == state; // @[Conditional.scala 37:30:@1094.10]
  assign _GEN_8 = io_done ? 2'h0 : 2'h2; // @[GunzipOutBuf.scala 75:22:@1096.12]
  assign _GEN_9 = _T_38 ? _GEN_8 : state; // @[Conditional.scala 39:67:@1095.10]
  assign _GEN_10 = _T_37 ? _GEN_7 : _GEN_9; // @[Conditional.scala 39:67:@1088.8]
  assign _GEN_11 = _T_36 ? 2'h2 : _GEN_10; // @[Conditional.scala 39:67:@1083.6]
  assign _GEN_12 = _T_35 ? _GEN_6 : _GEN_11; // @[Conditional.scala 40:58:@1076.4]
  assign _T_39 = state == 2'h0; // @[GunzipOutBuf.scala 83:15:@1103.4]
  assign _T_40 = _T_39 & io_enable; // @[GunzipOutBuf.scala 83:25:@1104.4]
  assign _T_41 = out_buf_wr_pos - io_dist; // @[GunzipOutBuf.scala 84:38:@1106.6]
  assign _T_42 = $unsigned(_T_41); // @[GunzipOutBuf.scala 84:38:@1107.6]
  assign _T_43 = _T_42[14:0]; // @[GunzipOutBuf.scala 84:38:@1108.6]
  assign _T_44 = state == 2'h2; // @[GunzipOutBuf.scala 86:22:@1113.6]
  assign _T_45 = _T_44 & io_data_out_ready; // @[GunzipOutBuf.scala 86:32:@1114.6]
  assign _T_47 = out_buf_rd_pos + 15'h1; // @[GunzipOutBuf.scala 87:38:@1116.8]
  assign _T_48 = out_buf_rd_pos + 15'h1; // @[GunzipOutBuf.scala 87:38:@1117.8]
  assign _T_50 = rem_len - 15'h1; // @[GunzipOutBuf.scala 88:24:@1119.8]
  assign _T_51 = $unsigned(_T_50); // @[GunzipOutBuf.scala 88:24:@1120.8]
  assign _T_52 = _T_51[14:0]; // @[GunzipOutBuf.scala 88:24:@1121.8]
  assign _GEN_13 = _T_45 ? _T_48 : out_buf_rd_pos; // @[GunzipOutBuf.scala 86:54:@1115.6]
  assign _GEN_14 = _T_45 ? _T_52 : rem_len; // @[GunzipOutBuf.scala 86:54:@1115.6]
  assign _GEN_15 = _T_40 ? _T_43 : _GEN_13; // @[GunzipOutBuf.scala 83:39:@1105.4]
  assign _T_61 = state == 2'h3; // @[GunzipOutBuf.scala 94:20:@1135.4]
  assign _T_63 = rem_len == 15'h0; // @[GunzipOutBuf.scala 94:42:@1136.4]
  assign io_done = _T_61 & _T_63; // @[GunzipOutBuf.scala 94:11:@1138.4]
  assign io_data_out_bits = out_buf__T_59_data; // @[GunzipOutBuf.scala 91:20:@1132.4]
  assign io_data_out_valid = state == 2'h2; // @[GunzipOutBuf.scala 92:21:@1134.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32768; initvar = initvar+1)
    out_buf[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  out_buf_wr_pos = _RAND_1[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_buf_rd_pos = _RAND_2[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  rem_len = _RAND_3[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_buf__T_59_addr_pipe_0 = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(out_buf__T_30_en & out_buf__T_30_mask) begin
      out_buf[out_buf__T_30_addr] <= out_buf__T_30_data; // @[GunzipOutBuf.scala 46:28:@1063.4]
    end
    if (reset) begin
      out_buf_wr_pos <= 15'h0;
    end else begin
      if (io_valid_in) begin
        out_buf_wr_pos <= _T_33;
      end
    end
    if (reset) begin
      out_buf_rd_pos <= 15'h0;
    end else begin
      if (_T_40) begin
        out_buf_rd_pos <= _T_43;
      end else begin
        if (_T_45) begin
          out_buf_rd_pos <= _T_48;
        end
      end
    end
    if (_T_40) begin
      rem_len <= io_len;
    end else begin
      if (_T_45) begin
        rem_len <= _T_52;
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_35) begin
        if (io_enable) begin
          state <= 2'h1;
        end
      end else begin
        if (_T_36) begin
          state <= 2'h2;
        end else begin
          if (_T_37) begin
            if (io_data_out_ready) begin
              state <= 2'h3;
            end
          end else begin
            if (_T_38) begin
              if (io_done) begin
                state <= 2'h0;
              end else begin
                state <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (_GEN_3) begin
      out_buf__T_59_addr_pipe_0 <= out_buf_rd_pos;
    end
  end
endmodule
module GunzipEngine( // @[:@1140.2]
  input        clock, // @[:@1141.4]
  input        reset, // @[:@1142.4]
  output       io_data_in_ready, // @[:@1143.4]
  input        io_data_in_valid, // @[:@1143.4]
  input  [7:0] io_data_in_bits, // @[:@1143.4]
  input        io_data_out_ready, // @[:@1143.4]
  output       io_data_out_valid, // @[:@1143.4]
  output [7:0] io_data_out_bits_data, // @[:@1143.4]
  output       io_data_out_bits_last // @[:@1143.4]
);
  wire  bit_skipper_clock; // @[GunzipEngine.scala 45:27:@1208.4]
  wire  bit_skipper_reset; // @[GunzipEngine.scala 45:27:@1208.4]
  wire  bit_skipper_io_data_in_valid; // @[GunzipEngine.scala 45:27:@1208.4]
  wire  bit_skipper_io_data_in_ready; // @[GunzipEngine.scala 45:27:@1208.4]
  wire  bit_skipper_io_done; // @[GunzipEngine.scala 45:27:@1208.4]
  wire  dec_lit_clock; // @[GunzipEngine.scala 52:23:@1213.4]
  wire  dec_lit_reset; // @[GunzipEngine.scala 52:23:@1213.4]
  wire  dec_lit_io_data_in_valid; // @[GunzipEngine.scala 52:23:@1213.4]
  wire  dec_lit_io_data_in_ready; // @[GunzipEngine.scala 52:23:@1213.4]
  wire  dec_lit_io_data_in_bits; // @[GunzipEngine.scala 52:23:@1213.4]
  wire  dec_lit_io_enable; // @[GunzipEngine.scala 52:23:@1213.4]
  wire [8:0] dec_lit_io_data; // @[GunzipEngine.scala 52:23:@1213.4]
  wire  dec_lit_io_valid; // @[GunzipEngine.scala 52:23:@1213.4]
  wire  lut_len_clock; // @[GunzipEngine.scala 66:23:@1221.4]
  wire  lut_len_reset; // @[GunzipEngine.scala 66:23:@1221.4]
  wire  lut_len_io_data_in_valid; // @[GunzipEngine.scala 66:23:@1221.4]
  wire  lut_len_io_data_in_ready; // @[GunzipEngine.scala 66:23:@1221.4]
  wire  lut_len_io_data_in_bits; // @[GunzipEngine.scala 66:23:@1221.4]
  wire  lut_len_io_enable; // @[GunzipEngine.scala 66:23:@1221.4]
  wire [8:0] lut_len_io_lut_idx; // @[GunzipEngine.scala 66:23:@1221.4]
  wire  lut_len_io_done; // @[GunzipEngine.scala 66:23:@1221.4]
  wire [14:0] lut_len_io_lut_out; // @[GunzipEngine.scala 66:23:@1221.4]
  wire  dec_dist_clock; // @[GunzipEngine.scala 76:24:@1233.4]
  wire  dec_dist_reset; // @[GunzipEngine.scala 76:24:@1233.4]
  wire  dec_dist_io_data_in_valid; // @[GunzipEngine.scala 76:24:@1233.4]
  wire  dec_dist_io_data_in_ready; // @[GunzipEngine.scala 76:24:@1233.4]
  wire  dec_dist_io_data_in_bits; // @[GunzipEngine.scala 76:24:@1233.4]
  wire  dec_dist_io_enable; // @[GunzipEngine.scala 76:24:@1233.4]
  wire [8:0] dec_dist_io_data; // @[GunzipEngine.scala 76:24:@1233.4]
  wire  dec_dist_io_valid; // @[GunzipEngine.scala 76:24:@1233.4]
  wire  lut_dist_clock; // @[GunzipEngine.scala 91:24:@1241.4]
  wire  lut_dist_reset; // @[GunzipEngine.scala 91:24:@1241.4]
  wire  lut_dist_io_data_in_valid; // @[GunzipEngine.scala 91:24:@1241.4]
  wire  lut_dist_io_data_in_ready; // @[GunzipEngine.scala 91:24:@1241.4]
  wire  lut_dist_io_data_in_bits; // @[GunzipEngine.scala 91:24:@1241.4]
  wire  lut_dist_io_enable; // @[GunzipEngine.scala 91:24:@1241.4]
  wire [8:0] lut_dist_io_lut_idx; // @[GunzipEngine.scala 91:24:@1241.4]
  wire  lut_dist_io_done; // @[GunzipEngine.scala 91:24:@1241.4]
  wire [14:0] lut_dist_io_lut_out; // @[GunzipEngine.scala 91:24:@1241.4]
  wire  out_buf_clock; // @[GunzipEngine.scala 99:23:@1249.4]
  wire  out_buf_reset; // @[GunzipEngine.scala 99:23:@1249.4]
  wire [7:0] out_buf_io_data_in; // @[GunzipEngine.scala 99:23:@1249.4]
  wire  out_buf_io_valid_in; // @[GunzipEngine.scala 99:23:@1249.4]
  wire [14:0] out_buf_io_dist; // @[GunzipEngine.scala 99:23:@1249.4]
  wire [14:0] out_buf_io_len; // @[GunzipEngine.scala 99:23:@1249.4]
  wire  out_buf_io_enable; // @[GunzipEngine.scala 99:23:@1249.4]
  wire  out_buf_io_done; // @[GunzipEngine.scala 99:23:@1249.4]
  wire [7:0] out_buf_io_data_out_bits; // @[GunzipEngine.scala 99:23:@1249.4]
  wire  out_buf_io_data_out_valid; // @[GunzipEngine.scala 99:23:@1249.4]
  wire  out_buf_io_data_out_ready; // @[GunzipEngine.scala 99:23:@1249.4]
  wire [9:0] _T_126; // @[GunzipEngine.scala 70:41:@1228.4]
  wire [9:0] _T_127; // @[GunzipEngine.scala 70:41:@1229.4]
  reg [2:0] state; // @[GunzipEngine.scala 112:22:@1259.4]
  reg [31:0] _RAND_0;
  reg [7:0] out_data; // @[GunzipEngine.scala 114:21:@1260.4]
  reg [31:0] _RAND_1;
  reg  out_valid; // @[GunzipEngine.scala 115:22:@1261.4]
  reg [31:0] _RAND_2;
  reg  out_last; // @[GunzipEngine.scala 116:21:@1262.4]
  reg [31:0] _RAND_3;
  wire  _T_146; // @[Conditional.scala 37:30:@1270.4]
  wire  _T_149; // @[GunzipEngine.scala 130:15:@1275.8]
  wire [2:0] _GEN_0; // @[GunzipEngine.scala 128:34:@1272.6]
  wire  _T_150; // @[Conditional.scala 37:30:@1282.6]
  wire  _T_153; // @[GunzipEngine.scala 136:31:@1286.10]
  wire [7:0] _T_154; // @[GunzipEngine.scala 137:38:@1288.12]
  wire  _T_157; // @[GunzipEngine.scala 139:38:@1293.12]
  wire [2:0] _GEN_3; // @[GunzipEngine.scala 139:49:@1294.12]
  wire [7:0] _GEN_4; // @[GunzipEngine.scala 136:40:@1287.10]
  wire  _GEN_5; // @[GunzipEngine.scala 136:40:@1287.10]
  wire  _GEN_6; // @[GunzipEngine.scala 136:40:@1287.10]
  wire [2:0] _GEN_7; // @[GunzipEngine.scala 136:40:@1287.10]
  wire [7:0] _GEN_8; // @[GunzipEngine.scala 135:31:@1285.8]
  wire  _GEN_9; // @[GunzipEngine.scala 135:31:@1285.8]
  wire  _GEN_10; // @[GunzipEngine.scala 135:31:@1285.8]
  wire [2:0] _GEN_11; // @[GunzipEngine.scala 135:31:@1285.8]
  wire  _T_161; // @[Conditional.scala 37:30:@1305.8]
  wire [2:0] _GEN_12; // @[GunzipEngine.scala 150:30:@1308.10]
  wire  _T_166; // @[Conditional.scala 37:30:@1318.10]
  wire [2:0] _GEN_13; // @[GunzipEngine.scala 157:32:@1321.12]
  wire  _T_168; // @[Conditional.scala 37:30:@1326.12]
  wire [2:0] _GEN_14; // @[GunzipEngine.scala 163:31:@1329.14]
  wire  _T_173; // @[Conditional.scala 37:30:@1339.14]
  wire [2:0] _GEN_15; // @[GunzipEngine.scala 173:30:@1344.16]
  wire  _GEN_17; // @[Conditional.scala 39:67:@1340.14]
  wire [7:0] _GEN_18; // @[Conditional.scala 39:67:@1340.14]
  wire [2:0] _GEN_19; // @[Conditional.scala 39:67:@1340.14]
  wire [2:0] _GEN_21; // @[Conditional.scala 39:67:@1327.12]
  wire  _GEN_22; // @[Conditional.scala 39:67:@1327.12]
  wire  _GEN_23; // @[Conditional.scala 39:67:@1327.12]
  wire [7:0] _GEN_24; // @[Conditional.scala 39:67:@1327.12]
  wire [2:0] _GEN_26; // @[Conditional.scala 39:67:@1319.10]
  wire  _GEN_27; // @[Conditional.scala 39:67:@1319.10]
  wire  _GEN_28; // @[Conditional.scala 39:67:@1319.10]
  wire  _GEN_29; // @[Conditional.scala 39:67:@1319.10]
  wire [7:0] _GEN_30; // @[Conditional.scala 39:67:@1319.10]
  wire [2:0] _GEN_32; // @[Conditional.scala 39:67:@1306.8]
  wire  _GEN_33; // @[Conditional.scala 39:67:@1306.8]
  wire  _GEN_34; // @[Conditional.scala 39:67:@1306.8]
  wire  _GEN_35; // @[Conditional.scala 39:67:@1306.8]
  wire  _GEN_36; // @[Conditional.scala 39:67:@1306.8]
  wire [7:0] _GEN_37; // @[Conditional.scala 39:67:@1306.8]
  wire [7:0] _GEN_39; // @[Conditional.scala 39:67:@1283.6]
  wire  _GEN_40; // @[Conditional.scala 39:67:@1283.6]
  wire  _GEN_41; // @[Conditional.scala 39:67:@1283.6]
  wire [2:0] _GEN_42; // @[Conditional.scala 39:67:@1283.6]
  wire  _GEN_43; // @[Conditional.scala 39:67:@1283.6]
  wire  _GEN_44; // @[Conditional.scala 39:67:@1283.6]
  wire  _GEN_45; // @[Conditional.scala 39:67:@1283.6]
  wire  _GEN_46; // @[Conditional.scala 39:67:@1283.6]
  wire [2:0] _GEN_47; // @[Conditional.scala 40:58:@1271.4]
  wire  _T_176; // @[GunzipEngine.scala 184:15:@1352.4]
  wire  _GEN_56; // @[GunzipEngine.scala 184:26:@1353.4]
  wire  _T_177; // @[GunzipEngine.scala 187:15:@1356.4]
  wire  _GEN_57; // @[GunzipEngine.scala 187:28:@1357.4]
  wire  _T_178; // @[GunzipEngine.scala 190:15:@1360.4]
  wire  _GEN_58; // @[GunzipEngine.scala 190:25:@1361.4]
  wire  _T_179; // @[GunzipEngine.scala 193:15:@1364.4]
  wire  _GEN_59; // @[GunzipEngine.scala 193:29:@1365.4]
  wire  _T_180; // @[GunzipEngine.scala 196:15:@1368.4]
  wire  _GEN_61; // @[GunzipEngine.scala 130:15:@1277.10]
  wire  _GEN_62; // @[GunzipEngine.scala 152:15:@1313.14]
  wire  _GEN_63; // @[GunzipEngine.scala 152:15:@1313.14]
  wire  _GEN_64; // @[GunzipEngine.scala 152:15:@1313.14]
  wire  _GEN_65; // @[GunzipEngine.scala 152:15:@1313.14]
  wire  _GEN_66; // @[GunzipEngine.scala 152:15:@1313.14]
  wire  _GEN_70; // @[GunzipEngine.scala 165:15:@1334.18]
  wire  _GEN_71; // @[GunzipEngine.scala 165:15:@1334.18]
  wire  _GEN_72; // @[GunzipEngine.scala 165:15:@1334.18]
  wire  _GEN_73; // @[GunzipEngine.scala 165:15:@1334.18]
  wire  _GEN_74; // @[GunzipEngine.scala 165:15:@1334.18]
  wire  _GEN_75; // @[GunzipEngine.scala 165:15:@1334.18]
  GunzipBitSkipper bit_skipper ( // @[GunzipEngine.scala 45:27:@1208.4]
    .clock(bit_skipper_clock),
    .reset(bit_skipper_reset),
    .io_data_in_valid(bit_skipper_io_data_in_valid),
    .io_data_in_ready(bit_skipper_io_data_in_ready),
    .io_done(bit_skipper_io_done)
  );
  GunzipHuffDecoder dec_lit ( // @[GunzipEngine.scala 52:23:@1213.4]
    .clock(dec_lit_clock),
    .reset(dec_lit_reset),
    .io_data_in_valid(dec_lit_io_data_in_valid),
    .io_data_in_ready(dec_lit_io_data_in_ready),
    .io_data_in_bits(dec_lit_io_data_in_bits),
    .io_enable(dec_lit_io_enable),
    .io_data(dec_lit_io_data),
    .io_valid(dec_lit_io_valid)
  );
  GunzipLenDistLut lut_len ( // @[GunzipEngine.scala 66:23:@1221.4]
    .clock(lut_len_clock),
    .reset(lut_len_reset),
    .io_data_in_valid(lut_len_io_data_in_valid),
    .io_data_in_ready(lut_len_io_data_in_ready),
    .io_data_in_bits(lut_len_io_data_in_bits),
    .io_enable(lut_len_io_enable),
    .io_lut_idx(lut_len_io_lut_idx),
    .io_done(lut_len_io_done),
    .io_lut_out(lut_len_io_lut_out)
  );
  GunzipHuffDecoder_1 dec_dist ( // @[GunzipEngine.scala 76:24:@1233.4]
    .clock(dec_dist_clock),
    .reset(dec_dist_reset),
    .io_data_in_valid(dec_dist_io_data_in_valid),
    .io_data_in_ready(dec_dist_io_data_in_ready),
    .io_data_in_bits(dec_dist_io_data_in_bits),
    .io_enable(dec_dist_io_enable),
    .io_data(dec_dist_io_data),
    .io_valid(dec_dist_io_valid)
  );
  GunzipLenDistLut_1 lut_dist ( // @[GunzipEngine.scala 91:24:@1241.4]
    .clock(lut_dist_clock),
    .reset(lut_dist_reset),
    .io_data_in_valid(lut_dist_io_data_in_valid),
    .io_data_in_ready(lut_dist_io_data_in_ready),
    .io_data_in_bits(lut_dist_io_data_in_bits),
    .io_enable(lut_dist_io_enable),
    .io_lut_idx(lut_dist_io_lut_idx),
    .io_done(lut_dist_io_done),
    .io_lut_out(lut_dist_io_lut_out)
  );
  GunzipOutBuf out_buf ( // @[GunzipEngine.scala 99:23:@1249.4]
    .clock(out_buf_clock),
    .reset(out_buf_reset),
    .io_data_in(out_buf_io_data_in),
    .io_valid_in(out_buf_io_valid_in),
    .io_dist(out_buf_io_dist),
    .io_len(out_buf_io_len),
    .io_enable(out_buf_io_enable),
    .io_done(out_buf_io_done),
    .io_data_out_bits(out_buf_io_data_out_bits),
    .io_data_out_valid(out_buf_io_data_out_valid),
    .io_data_out_ready(out_buf_io_data_out_ready)
  );
  assign _T_126 = dec_lit_io_data - 9'h101; // @[GunzipEngine.scala 70:41:@1228.4]
  assign _T_127 = $unsigned(_T_126); // @[GunzipEngine.scala 70:41:@1229.4]
  assign _T_146 = 3'h0 == state; // @[Conditional.scala 37:30:@1270.4]
  assign _T_149 = reset == 1'h0; // @[GunzipEngine.scala 130:15:@1275.8]
  assign _GEN_0 = bit_skipper_io_done ? 3'h1 : state; // @[GunzipEngine.scala 128:34:@1272.6]
  assign _T_150 = 3'h1 == state; // @[Conditional.scala 37:30:@1282.6]
  assign _T_153 = dec_lit_io_data < 9'h100; // @[GunzipEngine.scala 136:31:@1286.10]
  assign _T_154 = dec_lit_io_data[7:0]; // @[GunzipEngine.scala 137:38:@1288.12]
  assign _T_157 = dec_lit_io_data == 9'h100; // @[GunzipEngine.scala 139:38:@1293.12]
  assign _GEN_3 = _T_157 ? state : 3'h2; // @[GunzipEngine.scala 139:49:@1294.12]
  assign _GEN_4 = _T_153 ? _T_154 : 8'h0; // @[GunzipEngine.scala 136:40:@1287.10]
  assign _GEN_5 = _T_153 ? 1'h1 : _T_157; // @[GunzipEngine.scala 136:40:@1287.10]
  assign _GEN_6 = _T_153 ? 1'h0 : _T_157; // @[GunzipEngine.scala 136:40:@1287.10]
  assign _GEN_7 = _T_153 ? state : _GEN_3; // @[GunzipEngine.scala 136:40:@1287.10]
  assign _GEN_8 = dec_lit_io_valid ? _GEN_4 : 8'h0; // @[GunzipEngine.scala 135:31:@1285.8]
  assign _GEN_9 = dec_lit_io_valid ? _GEN_5 : 1'h0; // @[GunzipEngine.scala 135:31:@1285.8]
  assign _GEN_10 = dec_lit_io_valid ? _GEN_6 : 1'h0; // @[GunzipEngine.scala 135:31:@1285.8]
  assign _GEN_11 = dec_lit_io_valid ? _GEN_7 : state; // @[GunzipEngine.scala 135:31:@1285.8]
  assign _T_161 = 3'h2 == state; // @[Conditional.scala 37:30:@1305.8]
  assign _GEN_12 = lut_len_io_done ? 3'h3 : state; // @[GunzipEngine.scala 150:30:@1308.10]
  assign _T_166 = 3'h3 == state; // @[Conditional.scala 37:30:@1318.10]
  assign _GEN_13 = dec_dist_io_valid ? 3'h4 : state; // @[GunzipEngine.scala 157:32:@1321.12]
  assign _T_168 = 3'h4 == state; // @[Conditional.scala 37:30:@1326.12]
  assign _GEN_14 = lut_dist_io_done ? 3'h5 : state; // @[GunzipEngine.scala 163:31:@1329.14]
  assign _T_173 = 3'h5 == state; // @[Conditional.scala 37:30:@1339.14]
  assign _GEN_15 = out_buf_io_done ? 3'h1 : state; // @[GunzipEngine.scala 173:30:@1344.16]
  assign _GEN_17 = _T_173 ? out_buf_io_data_out_valid : 1'h0; // @[Conditional.scala 39:67:@1340.14]
  assign _GEN_18 = _T_173 ? out_buf_io_data_out_bits : 8'h0; // @[Conditional.scala 39:67:@1340.14]
  assign _GEN_19 = _T_173 ? _GEN_15 : state; // @[Conditional.scala 39:67:@1340.14]
  assign _GEN_21 = _T_168 ? _GEN_14 : _GEN_19; // @[Conditional.scala 39:67:@1327.12]
  assign _GEN_22 = _T_168 ? 1'h0 : _T_173; // @[Conditional.scala 39:67:@1327.12]
  assign _GEN_23 = _T_168 ? 1'h0 : _GEN_17; // @[Conditional.scala 39:67:@1327.12]
  assign _GEN_24 = _T_168 ? 8'h0 : _GEN_18; // @[Conditional.scala 39:67:@1327.12]
  assign _GEN_26 = _T_166 ? _GEN_13 : _GEN_21; // @[Conditional.scala 39:67:@1319.10]
  assign _GEN_27 = _T_166 ? 1'h0 : _T_168; // @[Conditional.scala 39:67:@1319.10]
  assign _GEN_28 = _T_166 ? 1'h0 : _GEN_22; // @[Conditional.scala 39:67:@1319.10]
  assign _GEN_29 = _T_166 ? 1'h0 : _GEN_23; // @[Conditional.scala 39:67:@1319.10]
  assign _GEN_30 = _T_166 ? 8'h0 : _GEN_24; // @[Conditional.scala 39:67:@1319.10]
  assign _GEN_32 = _T_161 ? _GEN_12 : _GEN_26; // @[Conditional.scala 39:67:@1306.8]
  assign _GEN_33 = _T_161 ? 1'h0 : _T_166; // @[Conditional.scala 39:67:@1306.8]
  assign _GEN_34 = _T_161 ? 1'h0 : _GEN_27; // @[Conditional.scala 39:67:@1306.8]
  assign _GEN_35 = _T_161 ? 1'h0 : _GEN_28; // @[Conditional.scala 39:67:@1306.8]
  assign _GEN_36 = _T_161 ? 1'h0 : _GEN_29; // @[Conditional.scala 39:67:@1306.8]
  assign _GEN_37 = _T_161 ? 8'h0 : _GEN_30; // @[Conditional.scala 39:67:@1306.8]
  assign _GEN_39 = _T_150 ? _GEN_8 : _GEN_37; // @[Conditional.scala 39:67:@1283.6]
  assign _GEN_40 = _T_150 ? _GEN_9 : _GEN_36; // @[Conditional.scala 39:67:@1283.6]
  assign _GEN_41 = _T_150 ? _GEN_10 : 1'h0; // @[Conditional.scala 39:67:@1283.6]
  assign _GEN_42 = _T_150 ? _GEN_11 : _GEN_32; // @[Conditional.scala 39:67:@1283.6]
  assign _GEN_43 = _T_150 ? 1'h0 : _T_161; // @[Conditional.scala 39:67:@1283.6]
  assign _GEN_44 = _T_150 ? 1'h0 : _GEN_33; // @[Conditional.scala 39:67:@1283.6]
  assign _GEN_45 = _T_150 ? 1'h0 : _GEN_34; // @[Conditional.scala 39:67:@1283.6]
  assign _GEN_46 = _T_150 ? 1'h0 : _GEN_35; // @[Conditional.scala 39:67:@1283.6]
  assign _GEN_47 = _T_146 ? _GEN_0 : _GEN_42; // @[Conditional.scala 40:58:@1271.4]
  assign _T_176 = state == 3'h0; // @[GunzipEngine.scala 184:15:@1352.4]
  assign _GEN_56 = _T_176 ? bit_skipper_io_data_in_ready : 1'h0; // @[GunzipEngine.scala 184:26:@1353.4]
  assign _T_177 = state == 3'h1; // @[GunzipEngine.scala 187:15:@1356.4]
  assign _GEN_57 = _T_177 ? dec_lit_io_data_in_ready : _GEN_56; // @[GunzipEngine.scala 187:28:@1357.4]
  assign _T_178 = state == 3'h2; // @[GunzipEngine.scala 190:15:@1360.4]
  assign _GEN_58 = _T_178 ? lut_len_io_data_in_ready : _GEN_57; // @[GunzipEngine.scala 190:25:@1361.4]
  assign _T_179 = state == 3'h3; // @[GunzipEngine.scala 193:15:@1364.4]
  assign _GEN_59 = _T_179 ? dec_dist_io_data_in_ready : _GEN_58; // @[GunzipEngine.scala 193:29:@1365.4]
  assign _T_180 = state == 3'h4; // @[GunzipEngine.scala 196:15:@1368.4]
  assign io_data_in_ready = _T_180 ? lut_dist_io_data_in_ready : _GEN_59; // @[GunzipEngine.scala 183:20:@1351.4 GunzipEngine.scala 185:22:@1354.6 GunzipEngine.scala 188:22:@1358.6 GunzipEngine.scala 191:22:@1362.6 GunzipEngine.scala 194:22:@1366.6 GunzipEngine.scala 197:22:@1370.6]
  assign io_data_out_valid = out_valid; // @[GunzipEngine.scala 179:21:@1348.4]
  assign io_data_out_bits_data = out_data; // @[GunzipEngine.scala 180:25:@1349.4]
  assign io_data_out_bits_last = out_last; // @[GunzipEngine.scala 181:25:@1350.4]
  assign bit_skipper_clock = clock; // @[:@1209.4]
  assign bit_skipper_reset = reset; // @[:@1210.4]
  assign bit_skipper_io_data_in_valid = io_data_in_valid; // @[GunzipEngine.scala 46:32:@1211.4]
  assign dec_lit_clock = clock; // @[:@1214.4]
  assign dec_lit_reset = reset; // @[:@1215.4]
  assign dec_lit_io_data_in_valid = io_data_in_valid; // @[GunzipEngine.scala 53:28:@1216.4]
  assign dec_lit_io_data_in_bits = io_data_in_bits[0]; // @[GunzipEngine.scala 54:27:@1218.4]
  assign dec_lit_io_enable = _T_146 ? 1'h0 : _T_150; // @[GunzipEngine.scala 55:21:@1219.4]
  assign lut_len_clock = clock; // @[:@1222.4]
  assign lut_len_reset = reset; // @[:@1223.4]
  assign lut_len_io_data_in_valid = io_data_in_valid; // @[GunzipEngine.scala 68:28:@1226.4]
  assign lut_len_io_data_in_bits = io_data_in_bits[0]; // @[GunzipEngine.scala 67:27:@1225.4]
  assign lut_len_io_enable = _T_146 ? 1'h0 : _GEN_43; // @[GunzipEngine.scala 69:21:@1227.4]
  assign lut_len_io_lut_idx = _T_127[8:0]; // @[GunzipEngine.scala 70:22:@1231.4]
  assign dec_dist_clock = clock; // @[:@1234.4]
  assign dec_dist_reset = reset; // @[:@1235.4]
  assign dec_dist_io_data_in_valid = io_data_in_valid; // @[GunzipEngine.scala 77:29:@1236.4]
  assign dec_dist_io_data_in_bits = io_data_in_bits[0]; // @[GunzipEngine.scala 78:28:@1238.4]
  assign dec_dist_io_enable = _T_146 ? 1'h0 : _GEN_44; // @[GunzipEngine.scala 79:22:@1239.4]
  assign lut_dist_clock = clock; // @[:@1242.4]
  assign lut_dist_reset = reset; // @[:@1243.4]
  assign lut_dist_io_data_in_valid = io_data_in_valid; // @[GunzipEngine.scala 93:29:@1246.4]
  assign lut_dist_io_data_in_bits = io_data_in_bits[0]; // @[GunzipEngine.scala 92:28:@1245.4]
  assign lut_dist_io_enable = _T_146 ? 1'h0 : _GEN_45; // @[GunzipEngine.scala 94:22:@1247.4]
  assign lut_dist_io_lut_idx = dec_dist_io_data; // @[GunzipEngine.scala 95:23:@1248.4]
  assign out_buf_clock = clock; // @[:@1250.4]
  assign out_buf_reset = reset; // @[:@1251.4]
  assign out_buf_io_data_in = io_data_out_bits_data; // @[GunzipEngine.scala 100:22:@1252.4]
  assign out_buf_io_valid_in = io_data_out_valid & io_data_out_ready; // @[GunzipEngine.scala 101:23:@1254.4]
  assign out_buf_io_dist = lut_dist_io_lut_out; // @[GunzipEngine.scala 103:19:@1255.4]
  assign out_buf_io_len = lut_len_io_lut_out; // @[GunzipEngine.scala 104:19:@1256.4]
  assign out_buf_io_enable = _T_146 ? 1'h0 : _GEN_46; // @[GunzipEngine.scala 105:21:@1257.4 GunzipEngine.scala 169:25:@1341.16]
  assign out_buf_io_data_out_ready = io_data_out_ready; // @[GunzipEngine.scala 107:29:@1258.4]
  assign _GEN_61 = _T_146 & bit_skipper_io_done; // @[GunzipEngine.scala 130:15:@1277.10]
  assign _GEN_62 = _T_146 == 1'h0; // @[GunzipEngine.scala 152:15:@1313.14]
  assign _GEN_63 = _T_150 == 1'h0; // @[GunzipEngine.scala 152:15:@1313.14]
  assign _GEN_64 = _GEN_62 & _GEN_63; // @[GunzipEngine.scala 152:15:@1313.14]
  assign _GEN_65 = _GEN_64 & _T_161; // @[GunzipEngine.scala 152:15:@1313.14]
  assign _GEN_66 = _GEN_65 & lut_len_io_done; // @[GunzipEngine.scala 152:15:@1313.14]
  assign _GEN_70 = _T_161 == 1'h0; // @[GunzipEngine.scala 165:15:@1334.18]
  assign _GEN_71 = _GEN_64 & _GEN_70; // @[GunzipEngine.scala 165:15:@1334.18]
  assign _GEN_72 = _T_166 == 1'h0; // @[GunzipEngine.scala 165:15:@1334.18]
  assign _GEN_73 = _GEN_71 & _GEN_72; // @[GunzipEngine.scala 165:15:@1334.18]
  assign _GEN_74 = _GEN_73 & _T_168; // @[GunzipEngine.scala 165:15:@1334.18]
  assign _GEN_75 = _GEN_74 & lut_dist_io_done; // @[GunzipEngine.scala 165:15:@1334.18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  out_data = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_valid = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_last = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      state <= 3'h0;
    end else begin
      if (_T_146) begin
        if (bit_skipper_io_done) begin
          state <= 3'h1;
        end
      end else begin
        if (_T_150) begin
          if (dec_lit_io_valid) begin
            if (!(_T_153)) begin
              if (!(_T_157)) begin
                state <= 3'h2;
              end
            end
          end
        end else begin
          if (_T_161) begin
            if (lut_len_io_done) begin
              state <= 3'h3;
            end
          end else begin
            if (_T_166) begin
              if (dec_dist_io_valid) begin
                state <= 3'h4;
              end
            end else begin
              if (_T_168) begin
                if (lut_dist_io_done) begin
                  state <= 3'h5;
                end
              end else begin
                if (_T_173) begin
                  if (out_buf_io_done) begin
                    state <= 3'h1;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_146) begin
      out_data <= 8'h0;
    end else begin
      if (_T_150) begin
        if (dec_lit_io_valid) begin
          if (_T_153) begin
            out_data <= _T_154;
          end else begin
            out_data <= 8'h0;
          end
        end else begin
          out_data <= 8'h0;
        end
      end else begin
        if (_T_161) begin
          out_data <= 8'h0;
        end else begin
          if (_T_166) begin
            out_data <= 8'h0;
          end else begin
            if (_T_168) begin
              out_data <= 8'h0;
            end else begin
              if (_T_173) begin
                out_data <= out_buf_io_data_out_bits;
              end else begin
                out_data <= 8'h0;
              end
            end
          end
        end
      end
    end
    if (_T_146) begin
      out_valid <= 1'h0;
    end else begin
      if (_T_150) begin
        if (dec_lit_io_valid) begin
          if (_T_153) begin
            out_valid <= 1'h1;
          end else begin
            out_valid <= _T_157;
          end
        end else begin
          out_valid <= 1'h0;
        end
      end else begin
        if (_T_161) begin
          out_valid <= 1'h0;
        end else begin
          if (_T_166) begin
            out_valid <= 1'h0;
          end else begin
            if (_T_168) begin
              out_valid <= 1'h0;
            end else begin
              if (_T_173) begin
                out_valid <= out_buf_io_data_out_valid;
              end else begin
                out_valid <= 1'h0;
              end
            end
          end
        end
      end
    end
    if (_T_146) begin
      out_last <= 1'h0;
    end else begin
      if (_T_150) begin
        if (dec_lit_io_valid) begin
          if (_T_153) begin
            out_last <= 1'h0;
          end else begin
            out_last <= _T_157;
          end
        end else begin
          out_last <= 1'h0;
        end
      end else begin
        out_last <= 1'h0;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_61 & _T_149) begin
          $fwrite(32'h80000002,"Bit skip finished\n"); // @[GunzipEngine.scala 130:15:@1277.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_66 & _T_149) begin
          $fwrite(32'h80000002,"  len: %d\n",lut_len_io_lut_out); // @[GunzipEngine.scala 152:15:@1313.14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_149) begin
          $fwrite(32'h80000002,"  dist: %d\n",lut_dist_io_lut_out); // @[GunzipEngine.scala 165:15:@1334.18]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
